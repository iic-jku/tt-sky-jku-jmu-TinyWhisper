* PEX produced on Sat Nov  8 09:20:06 PM CET 2025 using /foss/tools/sak/iic-pex.sh with m=1 and s=1
* NGSPICE file created from passive_voltage_mode_mixer.ext - technology: sky130A

.subckt passive_voltage_mode_mixer_pex vinp_IF VDD vinp_LO vinn_IF vout_RF VSS vinn_LO
X0 vinn_IF transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=23.12 ps=190.24001 w=1 l=0.15
X2 vout_RF transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=9.2 ps=74.4 w=1 l=0.15
X3 vout_RF transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X4 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=69.36 ps=478.23999 w=3 l=0.15
X5 transmission_gate_w_dummy_0.di_tg_ctrl lo_logic_0.inverter_NF6_0.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X6 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X7 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X8 vout_RF transmission_gate_w_dummy_2.di_tg_ctrl vinn_IF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X9 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X10 vout_RF transmission_gate_w_dummy_0.di_tg_ctrl_n vinp_IF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X11 vinp_IF transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X12 transmission_gate_w_dummy_0.di_tg_ctrl_n lo_logic_0.inverter_NF6_1.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X13 vout_RF transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=27.6 ps=186.39999 w=3 l=0.15
X14 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X15 transmission_gate_w_dummy_2.di_tg_ctrl lo_logic_1.inverter_NF6_0.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X16 vinn_IF transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X17 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X18 vout_RF transmission_gate_w_dummy_0.di_tg_ctrl vinp_IF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X19 VSS lo_logic_0.inv_cross lo_logic_0.inverter_NF6_1.vin VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X20 lo_logic_0.inverter_NF6_1.vin lo_logic_0.inv_cross VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X21 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X22 VDD lo_logic_1.transmission_gate_wo_dummy_0.v_b lo_logic_1.inv_cross VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X23 vinp_IF transmission_gate_w_dummy_0.di_tg_ctrl vinp_IF VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=13.8 ps=93.2 w=3 l=0.15
X24 transmission_gate_w_dummy_2.di_tg_ctrl_n lo_logic_1.inverter_NF6_1.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X25 lo_logic_0.inverter_NF6_0.vin lo_logic_0.buf_cross VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X26 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X27 vout_RF transmission_gate_w_dummy_0.di_tg_ctrl vinp_IF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X28 VDD lo_logic_1.inverter_NF6_1.vin transmission_gate_w_dummy_2.di_tg_ctrl_n VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X29 VDD lo_logic_0.inverter_NF6_1.vin transmission_gate_w_dummy_0.di_tg_ctrl_n VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X30 vout_RF transmission_gate_w_dummy_0.di_tg_ctrl_n vinp_IF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X31 vinp_IF transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X32 lo_logic_1.inverter_NF6_1.vin lo_logic_1.inv_cross VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X33 vout_RF transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X34 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X35 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X36 transmission_gate_w_dummy_0.di_tg_ctrl lo_logic_0.inverter_NF6_0.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X37 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X38 vinp_IF transmission_gate_w_dummy_0.di_tg_ctrl vinp_IF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X39 vinp_IF transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X40 VDD lo_logic_1.inverter_NF6_1.vin transmission_gate_w_dummy_2.di_tg_ctrl_n VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X41 VDD lo_logic_0.buf_cross lo_logic_0.inv_cross VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=3.81 ps=8.54 w=3 l=0.15
X42 transmission_gate_w_dummy_2.di_tg_ctrl_n lo_logic_1.inverter_NF6_1.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X43 transmission_gate_w_dummy_0.di_tg_ctrl lo_logic_0.inverter_NF6_0.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X44 lo_logic_0.transmission_gate_wo_dummy_0.v_b VSS vinp_LO VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.93 ps=6.62 w=3 l=0.15
X45 vinp_IF transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X46 vinp_IF transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X47 lo_logic_1.buf_cross lo_logic_1.inverter_NF2_1.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X48 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X49 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X50 VDD lo_logic_0.transmission_gate_wo_dummy_0.v_b lo_logic_0.inv_cross VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X51 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X52 vout_RF transmission_gate_w_dummy_0.di_tg_ctrl vinp_IF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X53 VDD lo_logic_0.inverter_NF6_0.vin transmission_gate_w_dummy_0.di_tg_ctrl VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X54 vout_RF transmission_gate_w_dummy_0.di_tg_ctrl_n vinp_IF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X55 vinp_IF transmission_gate_w_dummy_0.di_tg_ctrl_n vinp_IF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=4.6 ps=37.2 w=1 l=0.15
X56 VDD lo_logic_1.inv_cross lo_logic_1.inverter_NF6_1.vin VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X57 lo_logic_0.transmission_gate_wo_dummy_0.v_b VDD vinp_LO VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X58 lo_logic_1.buf_cross lo_logic_1.inverter_NF2_1.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X59 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X60 transmission_gate_w_dummy_2.di_tg_ctrl lo_logic_1.inverter_NF6_0.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X61 vinn_IF transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X62 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X63 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X64 vinn_IF transmission_gate_w_dummy_2.di_tg_ctrl vinn_IF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=13.8 ps=93.2 w=3 l=0.15
X65 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X66 VSS lo_logic_0.inverter_NF6_0.vin transmission_gate_w_dummy_0.di_tg_ctrl VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X67 vinp_LO VDD lo_logic_0.transmission_gate_wo_dummy_0.v_b VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X68 VSS lo_logic_1.inverter_NF6_1.vin transmission_gate_w_dummy_2.di_tg_ctrl_n VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X69 vout_RF transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X70 VSS lo_logic_1.inverter_NF6_0.vin transmission_gate_w_dummy_2.di_tg_ctrl VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X71 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X72 vout_RF transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X73 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X74 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X75 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X76 VSS lo_logic_0.buf_cross lo_logic_0.inv_cross VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=1.27 ps=4.54 w=1 l=0.15
X77 vout_RF transmission_gate_w_dummy_0.di_tg_ctrl vinp_IF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X78 vinn_IF transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X79 vinp_IF transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X80 VSS lo_logic_1.inverter_NF2_1.vin lo_logic_1.buf_cross VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X81 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X82 vinn_IF transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X83 VDD lo_logic_0.inv_cross lo_logic_0.inverter_NF6_1.vin VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X84 vinn_IF transmission_gate_w_dummy_2.di_tg_ctrl_n vinn_IF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=4.6 ps=37.2 w=1 l=0.15
X85 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X86 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X87 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X88 vout_RF transmission_gate_w_dummy_2.di_tg_ctrl_n vinn_IF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X89 vinp_IF transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X90 vout_RF transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X91 VDD lo_logic_1.inverter_NF2_1.vin lo_logic_1.buf_cross VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X92 transmission_gate_w_dummy_2.di_tg_ctrl lo_logic_1.inverter_NF6_0.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X93 VSS lo_logic_1.inverter_NF6_0.vin transmission_gate_w_dummy_2.di_tg_ctrl VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X94 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X95 VSS lo_logic_1.inv_cross lo_logic_1.buf_cross VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=1.27 ps=4.54 w=1 l=0.15
X96 vout_RF transmission_gate_w_dummy_2.di_tg_ctrl_n vinn_IF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X97 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X98 vinp_IF transmission_gate_w_dummy_0.di_tg_ctrl vinp_IF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X99 lo_logic_1.inverter_NF6_0.vin lo_logic_1.buf_cross VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X100 vinn_IF transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X101 vinn_IF transmission_gate_w_dummy_2.di_tg_ctrl vinn_IF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X102 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X103 vout_RF transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X104 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X105 VDD lo_logic_1.inverter_NF6_0.vin transmission_gate_w_dummy_2.di_tg_ctrl VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X106 transmission_gate_w_dummy_2.di_tg_ctrl_n lo_logic_1.inverter_NF6_1.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X107 vout_RF transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X108 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X109 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X110 vout_RF transmission_gate_w_dummy_2.di_tg_ctrl vinn_IF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X111 vout_RF transmission_gate_w_dummy_0.di_tg_ctrl vinp_IF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X112 vout_RF transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X113 vout_RF transmission_gate_w_dummy_2.di_tg_ctrl_n vinn_IF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X114 VSS lo_logic_0.inverter_NF6_1.vin transmission_gate_w_dummy_0.di_tg_ctrl_n VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X115 transmission_gate_w_dummy_0.di_tg_ctrl_n lo_logic_0.inverter_NF6_1.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X116 lo_logic_1.inverter_NF6_0.vin lo_logic_1.buf_cross VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X117 vout_RF transmission_gate_w_dummy_0.di_tg_ctrl_n vinp_IF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X118 vout_RF transmission_gate_w_dummy_2.di_tg_ctrl vinn_IF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X119 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X120 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X121 lo_logic_0.inv_cross lo_logic_0.transmission_gate_wo_dummy_0.v_b VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X122 transmission_gate_w_dummy_0.di_tg_ctrl_n lo_logic_0.inverter_NF6_1.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X123 VSS lo_logic_0.inverter_NF6_1.vin transmission_gate_w_dummy_0.di_tg_ctrl_n VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X124 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X125 vinn_IF transmission_gate_w_dummy_2.di_tg_ctrl_n vinn_IF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X126 vout_RF transmission_gate_w_dummy_2.di_tg_ctrl_n vinn_IF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X127 VDD vinp_LO lo_logic_0.inverter_NF2_1.vin VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X128 transmission_gate_w_dummy_0.di_tg_ctrl_n lo_logic_0.inverter_NF6_1.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X129 vinn_IF transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X130 transmission_gate_w_dummy_0.di_tg_ctrl lo_logic_0.inverter_NF6_0.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X131 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X132 vinp_IF transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X133 vinp_IF transmission_gate_w_dummy_0.di_tg_ctrl_n vinp_IF VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X134 VSS lo_logic_0.inverter_NF6_1.vin transmission_gate_w_dummy_0.di_tg_ctrl_n VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X135 vout_RF transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X136 vout_RF transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X137 vinn_IF transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X138 VDD lo_logic_1.inverter_NF6_0.vin transmission_gate_w_dummy_2.di_tg_ctrl VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X139 vout_RF transmission_gate_w_dummy_2.di_tg_ctrl vinn_IF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X140 VSS lo_logic_1.buf_cross lo_logic_1.inverter_NF6_0.vin VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X141 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X142 vout_RF transmission_gate_w_dummy_2.di_tg_ctrl vinn_IF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X143 vout_RF transmission_gate_w_dummy_0.di_tg_ctrl vinp_IF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X144 VSS lo_logic_0.inv_cross lo_logic_0.buf_cross VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=1.27 ps=4.54 w=1 l=0.15
X145 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X146 vinn_IF transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X147 VDD lo_logic_0.inverter_NF6_1.vin transmission_gate_w_dummy_0.di_tg_ctrl_n VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X148 vinp_IF transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X149 vout_RF transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X150 lo_logic_1.transmission_gate_wo_dummy_0.v_b VDD vinn_LO VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X151 vinn_IF transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X152 lo_logic_1.transmission_gate_wo_dummy_0.v_b VSS vinn_LO VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.93 ps=6.62 w=3 l=0.15
X153 vinp_IF transmission_gate_w_dummy_0.di_tg_ctrl_n vinp_IF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X154 VDD lo_logic_1.buf_cross lo_logic_1.inverter_NF6_0.vin VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X155 vinn_IF transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X156 VDD lo_logic_0.inverter_NF6_0.vin transmission_gate_w_dummy_0.di_tg_ctrl VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X157 vout_RF transmission_gate_w_dummy_0.di_tg_ctrl_n vinp_IF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X158 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X159 transmission_gate_w_dummy_2.di_tg_ctrl_n lo_logic_1.inverter_NF6_1.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X160 lo_logic_0.inverter_NF6_1.vin lo_logic_0.inv_cross VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X161 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X162 VSS vinp_LO lo_logic_0.inverter_NF2_1.vin VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X163 vout_RF transmission_gate_w_dummy_0.di_tg_ctrl_n vinp_IF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X164 vinp_IF transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X165 vinn_IF transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X166 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X167 transmission_gate_w_dummy_0.di_tg_ctrl_n lo_logic_0.inverter_NF6_1.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X168 vout_RF transmission_gate_w_dummy_0.di_tg_ctrl vinp_IF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X169 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X170 vout_RF transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X171 VDD lo_logic_0.inverter_NF2_1.vin lo_logic_0.buf_cross VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X172 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X173 VDD lo_logic_1.inverter_NF6_1.vin transmission_gate_w_dummy_2.di_tg_ctrl_n VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X174 vinp_IF transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X175 VDD lo_logic_1.inv_cross lo_logic_1.buf_cross VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=3.81 ps=8.54 w=3 l=0.15
X176 lo_logic_0.inverter_NF2_1.vin vinp_LO VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X177 VSS lo_logic_0.inverter_NF6_0.vin transmission_gate_w_dummy_0.di_tg_ctrl VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X178 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X179 lo_logic_1.inv_cross lo_logic_1.transmission_gate_wo_dummy_0.v_b VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X180 vout_RF transmission_gate_w_dummy_0.di_tg_ctrl_n vinp_IF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X181 vinp_IF transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X182 lo_logic_1.inverter_NF2_1.vin vinn_LO VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X183 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X184 vinp_LO VSS lo_logic_0.transmission_gate_wo_dummy_0.v_b VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0.495 ps=3.33 w=3 l=0.15
X185 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X186 transmission_gate_w_dummy_2.di_tg_ctrl lo_logic_1.inverter_NF6_0.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X187 transmission_gate_w_dummy_2.di_tg_ctrl_n lo_logic_1.inverter_NF6_1.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X188 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X189 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X190 vinp_IF transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X191 vinn_IF transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X192 transmission_gate_w_dummy_0.di_tg_ctrl_n lo_logic_0.inverter_NF6_1.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X193 vout_RF transmission_gate_w_dummy_0.di_tg_ctrl_n vinp_IF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X194 vout_RF transmission_gate_w_dummy_2.di_tg_ctrl_n vinn_IF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X195 VDD lo_logic_0.buf_cross lo_logic_0.inverter_NF6_0.vin VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X196 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X197 vinp_IF transmission_gate_w_dummy_0.di_tg_ctrl_n vinp_IF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X198 lo_logic_1.inverter_NF2_1.vin vinn_LO VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X199 VSS lo_logic_1.inverter_NF6_1.vin transmission_gate_w_dummy_2.di_tg_ctrl_n VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X200 transmission_gate_w_dummy_2.di_tg_ctrl_n lo_logic_1.inverter_NF6_1.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X201 VSS lo_logic_0.inverter_NF2_1.vin lo_logic_0.buf_cross VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X202 transmission_gate_w_dummy_0.di_tg_ctrl lo_logic_0.inverter_NF6_0.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X203 vinp_IF transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X204 VDD lo_logic_0.inv_cross lo_logic_0.buf_cross VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=3.81 ps=8.54 w=3 l=0.15
X205 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X206 VSS lo_logic_1.transmission_gate_wo_dummy_0.v_b lo_logic_1.inv_cross VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X207 lo_logic_0.inverter_NF2_1.vin vinp_LO VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X208 vinn_IF transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X209 vout_RF transmission_gate_w_dummy_2.di_tg_ctrl vinn_IF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X210 vinp_IF transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X211 vinn_IF transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X212 vinn_IF transmission_gate_w_dummy_2.di_tg_ctrl vinn_IF VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X213 vinp_IF transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X214 vout_RF transmission_gate_w_dummy_0.di_tg_ctrl vinp_IF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X215 VSS vinn_LO lo_logic_1.inverter_NF2_1.vin VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X216 VDD lo_logic_0.inverter_NF6_1.vin transmission_gate_w_dummy_0.di_tg_ctrl_n VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X217 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X218 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X219 VSS lo_logic_1.inverter_NF6_0.vin transmission_gate_w_dummy_2.di_tg_ctrl VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X220 VSS lo_logic_1.inverter_NF6_1.vin transmission_gate_w_dummy_2.di_tg_ctrl_n VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X221 vout_RF transmission_gate_w_dummy_2.di_tg_ctrl_n vinn_IF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X222 vout_RF transmission_gate_w_dummy_2.di_tg_ctrl_n vinn_IF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X223 vout_RF transmission_gate_w_dummy_0.di_tg_ctrl_n vinp_IF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X224 vinp_IF transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X225 transmission_gate_w_dummy_2.di_tg_ctrl lo_logic_1.inverter_NF6_0.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X226 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X227 lo_logic_1.inverter_NF6_1.vin lo_logic_1.inv_cross VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X228 lo_logic_0.buf_cross lo_logic_0.inverter_NF2_1.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X229 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X230 vinp_IF transmission_gate_w_dummy_0.di_tg_ctrl vinp_IF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X231 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X232 vinn_IF transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X233 VDD vinn_LO lo_logic_1.inverter_NF2_1.vin VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X234 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X235 vinn_IF transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X236 VSS lo_logic_0.buf_cross lo_logic_0.inverter_NF6_0.vin VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X237 vinn_LO VDD lo_logic_1.transmission_gate_wo_dummy_0.v_b VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X238 vinn_IF transmission_gate_w_dummy_2.di_tg_ctrl_n vinn_IF VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X239 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X240 vout_RF transmission_gate_w_dummy_2.di_tg_ctrl_n vinn_IF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X241 vinn_LO VSS lo_logic_1.transmission_gate_wo_dummy_0.v_b VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0.495 ps=3.33 w=3 l=0.15
X242 transmission_gate_w_dummy_0.di_tg_ctrl lo_logic_0.inverter_NF6_0.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X243 vinp_IF transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X244 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X245 vout_RF transmission_gate_w_dummy_2.di_tg_ctrl vinn_IF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X246 vout_RF transmission_gate_w_dummy_2.di_tg_ctrl vinn_IF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X247 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X248 VSS lo_logic_1.buf_cross lo_logic_1.inv_cross VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=1.27 ps=4.54 w=1 l=0.15
X249 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X250 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X251 vinn_IF transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X252 vout_RF transmission_gate_w_dummy_2.di_tg_ctrl_n vinn_IF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X253 vout_RF transmission_gate_w_dummy_0.di_tg_ctrl vinp_IF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X254 vinn_IF transmission_gate_w_dummy_2.di_tg_ctrl vinn_IF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X255 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X256 vout_RF transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X257 VDD lo_logic_0.inverter_NF6_0.vin transmission_gate_w_dummy_0.di_tg_ctrl VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X258 transmission_gate_w_dummy_2.di_tg_ctrl lo_logic_1.inverter_NF6_0.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X259 vout_RF transmission_gate_w_dummy_0.di_tg_ctrl_n vinp_IF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X260 VDD lo_logic_1.inverter_NF6_0.vin transmission_gate_w_dummy_2.di_tg_ctrl VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X261 vout_RF transmission_gate_w_dummy_2.di_tg_ctrl vinn_IF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X262 vout_RF transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X263 VDD lo_logic_1.buf_cross lo_logic_1.inv_cross VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=3.81 ps=8.54 w=3 l=0.15
X264 VSS lo_logic_1.inv_cross lo_logic_1.inverter_NF6_1.vin VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X265 vout_RF transmission_gate_w_dummy_0.di_tg_ctrl vinp_IF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X266 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X267 vout_RF transmission_gate_w_dummy_2.di_tg_ctrl_n vinn_IF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X268 lo_logic_0.inverter_NF6_0.vin lo_logic_0.buf_cross VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X269 vout_RF transmission_gate_w_dummy_2.di_tg_ctrl vinn_IF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X270 lo_logic_1.inv_cross lo_logic_1.transmission_gate_wo_dummy_0.v_b VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X271 VSS lo_logic_0.transmission_gate_wo_dummy_0.v_b lo_logic_0.inv_cross VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X272 lo_logic_0.buf_cross lo_logic_0.inverter_NF2_1.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X273 VSS lo_logic_0.inverter_NF6_0.vin transmission_gate_w_dummy_0.di_tg_ctrl VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X274 lo_logic_0.inv_cross lo_logic_0.transmission_gate_wo_dummy_0.v_b VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X275 vinn_IF transmission_gate_w_dummy_2.di_tg_ctrl_n vinn_IF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
C0 vinn_IF VSS 14.4924f
C1 vinn_LO VSS 4.18304f
C2 vout_RF VSS 30.7033f
C3 vinp_IF VSS 14.7225f
C4 vinp_LO VSS 4.18304f
C5 VDD VSS 0.19185p
C6 transmission_gate_w_dummy_2.di_tg_ctrl_n VSS 11.5065f
C7 lo_logic_1.inverter_NF6_1.vin VSS 4.48926f
C8 lo_logic_1.transmission_gate_wo_dummy_0.v_b VSS 2.83622f
C9 transmission_gate_w_dummy_2.di_tg_ctrl VSS 14.3155f
C10 lo_logic_1.inverter_NF6_0.vin VSS 4.48926f
C11 lo_logic_1.inv_cross VSS 7.66312f
C12 lo_logic_1.buf_cross VSS 7.89561f
C13 lo_logic_1.inverter_NF2_1.vin VSS 2.82434f
C14 transmission_gate_w_dummy_0.di_tg_ctrl_n VSS 11.5086f
C15 lo_logic_0.inverter_NF6_1.vin VSS 4.48926f
C16 lo_logic_0.transmission_gate_wo_dummy_0.v_b VSS 2.83622f
C17 transmission_gate_w_dummy_0.di_tg_ctrl VSS 14.3155f
C18 lo_logic_0.inverter_NF6_0.vin VSS 4.48926f
C19 lo_logic_0.inv_cross VSS 7.66312f
C20 lo_logic_0.buf_cross VSS 7.89561f
C21 lo_logic_0.inverter_NF2_1.vin VSS 2.82434f
.ends

