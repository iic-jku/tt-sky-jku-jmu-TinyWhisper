VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_TinyWhisper
  CLASS BLOCK ;
  FOREIGN tt_um_TinyWhisper ;
  ORIGIN 0.000 0.000 ;
  SIZE 334.880 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 73.599998 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.200000 ;
    ANTENNADIFFAREA 2.480000 ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.200000 ;
    ANTENNADIFFAREA 2.480000 ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.200000 ;
    ANTENNADIFFAREA 2.480000 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.200000 ;
    ANTENNADIFFAREA 2.480000 ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 96.000000 ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 231.050 158.995 254.950 159.000 ;
      LAYER pwell ;
        RECT 96.950 150.400 212.670 158.220 ;
      LAYER nwell ;
        RECT 231.050 153.805 254.960 158.995 ;
        RECT 231.050 153.800 254.950 153.805 ;
      LAYER pwell ;
        RECT 231.055 150.450 234.645 153.550 ;
        RECT 235.655 150.450 239.245 153.550 ;
        RECT 240.255 150.450 243.845 153.550 ;
        RECT 244.855 150.450 248.445 153.550 ;
        RECT 249.450 150.450 254.960 153.550 ;
      LAYER nwell ;
        RECT 231.050 149.695 254.950 149.700 ;
        RECT 75.280 136.720 84.690 147.910 ;
        RECT 86.030 136.720 98.020 147.910 ;
        RECT 99.355 136.720 111.345 147.910 ;
        RECT 112.680 136.720 122.090 147.910 ;
        RECT 123.430 136.720 135.420 147.910 ;
        RECT 136.755 136.720 148.745 147.910 ;
        RECT 150.080 136.720 162.070 147.910 ;
        RECT 163.405 136.720 175.395 147.910 ;
        RECT 176.730 136.720 188.720 147.910 ;
        RECT 190.055 136.720 199.465 147.910 ;
        RECT 200.805 136.720 212.795 147.910 ;
        RECT 214.130 136.720 226.120 147.910 ;
        RECT 231.050 144.505 254.960 149.695 ;
        RECT 256.625 148.100 271.255 153.290 ;
      LAYER pwell ;
        RECT 256.625 144.750 271.255 147.850 ;
      LAYER nwell ;
        RECT 231.050 144.500 254.950 144.505 ;
      LAYER pwell ;
        RECT 231.060 141.150 233.690 144.250 ;
        RECT 235.655 141.150 239.245 144.250 ;
        RECT 240.255 141.150 243.845 144.250 ;
        RECT 244.855 141.150 248.445 144.250 ;
        RECT 249.450 141.150 254.960 144.250 ;
      LAYER nwell ;
        RECT 231.050 138.145 254.950 138.150 ;
      LAYER pwell ;
        RECT 75.280 131.420 84.690 136.520 ;
        RECT 86.030 131.420 98.020 136.520 ;
        RECT 99.355 131.420 111.345 136.520 ;
        RECT 112.680 131.420 122.090 136.520 ;
        RECT 123.430 131.420 135.420 136.520 ;
        RECT 136.755 131.420 148.745 136.520 ;
        RECT 150.080 131.420 162.070 136.520 ;
        RECT 163.405 131.420 175.395 136.520 ;
        RECT 176.730 131.420 188.720 136.520 ;
        RECT 190.055 131.420 199.465 136.520 ;
        RECT 200.805 131.420 212.795 136.520 ;
        RECT 214.130 131.420 226.120 136.520 ;
      LAYER nwell ;
        RECT 231.050 132.955 254.960 138.145 ;
        RECT 231.050 132.950 254.950 132.955 ;
      LAYER pwell ;
        RECT 231.055 129.600 234.645 132.700 ;
        RECT 235.655 129.600 239.245 132.700 ;
        RECT 240.255 129.600 243.845 132.700 ;
        RECT 244.855 129.600 248.445 132.700 ;
        RECT 249.450 129.600 254.960 132.700 ;
        RECT 96.950 121.175 212.670 128.995 ;
      LAYER nwell ;
        RECT 231.050 128.845 254.950 128.850 ;
        RECT 231.050 123.655 254.960 128.845 ;
        RECT 256.625 127.250 271.255 132.440 ;
      LAYER pwell ;
        RECT 256.625 123.900 271.255 127.000 ;
      LAYER nwell ;
        RECT 231.050 123.650 254.950 123.655 ;
      LAYER pwell ;
        RECT 231.060 120.300 233.690 123.400 ;
        RECT 235.655 120.300 239.245 123.400 ;
        RECT 240.255 120.300 243.845 123.400 ;
        RECT 244.855 120.300 248.445 123.400 ;
        RECT 249.450 120.300 254.960 123.400 ;
      LAYER nwell ;
        RECT 231.050 105.495 254.950 105.500 ;
      LAYER pwell ;
        RECT 96.950 96.900 212.670 104.720 ;
      LAYER nwell ;
        RECT 231.050 100.305 254.960 105.495 ;
        RECT 231.050 100.300 254.950 100.305 ;
      LAYER pwell ;
        RECT 231.055 96.950 234.645 100.050 ;
        RECT 235.655 96.950 239.245 100.050 ;
        RECT 240.255 96.950 243.845 100.050 ;
        RECT 244.855 96.950 248.445 100.050 ;
        RECT 249.450 96.950 254.960 100.050 ;
      LAYER nwell ;
        RECT 231.050 96.195 254.950 96.200 ;
        RECT 75.280 83.220 84.690 94.410 ;
        RECT 86.030 83.220 98.020 94.410 ;
        RECT 99.355 83.220 111.345 94.410 ;
        RECT 112.680 83.220 122.090 94.410 ;
        RECT 123.430 83.220 135.420 94.410 ;
        RECT 136.755 83.220 148.745 94.410 ;
        RECT 150.080 83.220 162.070 94.410 ;
        RECT 163.405 83.220 175.395 94.410 ;
        RECT 176.730 83.220 188.720 94.410 ;
        RECT 190.055 83.220 199.465 94.410 ;
        RECT 200.805 83.220 212.795 94.410 ;
        RECT 214.130 83.220 226.120 94.410 ;
        RECT 231.050 91.005 254.960 96.195 ;
        RECT 256.625 94.600 271.255 99.790 ;
      LAYER pwell ;
        RECT 256.625 91.250 271.255 94.350 ;
      LAYER nwell ;
        RECT 231.050 91.000 254.950 91.005 ;
      LAYER pwell ;
        RECT 231.060 87.650 233.690 90.750 ;
        RECT 235.655 87.650 239.245 90.750 ;
        RECT 240.255 87.650 243.845 90.750 ;
        RECT 244.855 87.650 248.445 90.750 ;
        RECT 249.450 87.650 254.960 90.750 ;
      LAYER nwell ;
        RECT 231.050 84.645 254.950 84.650 ;
      LAYER pwell ;
        RECT 75.280 77.920 84.690 83.020 ;
        RECT 86.030 77.920 98.020 83.020 ;
        RECT 99.355 77.920 111.345 83.020 ;
        RECT 112.680 77.920 122.090 83.020 ;
        RECT 123.430 77.920 135.420 83.020 ;
        RECT 136.755 77.920 148.745 83.020 ;
        RECT 150.080 77.920 162.070 83.020 ;
        RECT 163.405 77.920 175.395 83.020 ;
        RECT 176.730 77.920 188.720 83.020 ;
        RECT 190.055 77.920 199.465 83.020 ;
        RECT 200.805 77.920 212.795 83.020 ;
        RECT 214.130 77.920 226.120 83.020 ;
      LAYER nwell ;
        RECT 231.050 79.455 254.960 84.645 ;
        RECT 231.050 79.450 254.950 79.455 ;
      LAYER pwell ;
        RECT 231.055 76.100 234.645 79.200 ;
        RECT 235.655 76.100 239.245 79.200 ;
        RECT 240.255 76.100 243.845 79.200 ;
        RECT 244.855 76.100 248.445 79.200 ;
        RECT 249.450 76.100 254.960 79.200 ;
        RECT 96.950 67.675 212.670 75.495 ;
      LAYER nwell ;
        RECT 231.050 75.345 254.950 75.350 ;
        RECT 231.050 70.155 254.960 75.345 ;
        RECT 256.625 73.750 271.255 78.940 ;
      LAYER pwell ;
        RECT 256.625 70.400 271.255 73.500 ;
      LAYER nwell ;
        RECT 231.050 70.150 254.950 70.155 ;
      LAYER pwell ;
        RECT 231.060 66.800 233.690 69.900 ;
        RECT 235.655 66.800 239.245 69.900 ;
        RECT 240.255 66.800 243.845 69.900 ;
        RECT 244.855 66.800 248.445 69.900 ;
        RECT 249.450 66.800 254.960 69.900 ;
      LAYER li1 ;
        RECT 75.275 157.870 228.050 159.850 ;
        RECT 231.050 158.995 271.250 159.850 ;
        RECT 75.275 150.750 97.300 157.870 ;
        RECT 97.780 155.230 98.130 157.390 ;
        RECT 98.610 155.230 98.960 157.390 ;
        RECT 99.440 155.230 99.790 157.390 ;
        RECT 100.270 155.230 100.620 157.390 ;
        RECT 101.100 155.230 101.450 157.390 ;
        RECT 101.930 155.230 102.280 157.390 ;
        RECT 102.760 155.230 103.110 157.390 ;
        RECT 103.590 155.230 103.940 157.390 ;
        RECT 104.420 155.230 104.770 157.390 ;
        RECT 105.250 155.230 105.600 157.390 ;
        RECT 106.080 155.230 106.430 157.390 ;
        RECT 106.910 155.230 107.260 157.390 ;
        RECT 107.740 155.230 108.090 157.390 ;
        RECT 108.570 155.230 108.920 157.390 ;
        RECT 109.400 155.230 109.750 157.390 ;
        RECT 110.230 155.230 110.580 157.390 ;
        RECT 111.060 155.230 111.410 157.390 ;
        RECT 111.890 155.230 112.240 157.390 ;
        RECT 112.720 155.230 113.070 157.390 ;
        RECT 113.550 155.230 113.900 157.390 ;
        RECT 114.380 155.230 114.730 157.390 ;
        RECT 115.210 155.230 115.560 157.390 ;
        RECT 116.040 155.230 116.390 157.390 ;
        RECT 116.870 155.230 117.220 157.390 ;
        RECT 117.700 155.230 118.050 157.390 ;
        RECT 118.530 155.230 118.880 157.390 ;
        RECT 119.360 155.230 119.710 157.390 ;
        RECT 120.190 155.230 120.540 157.390 ;
        RECT 121.020 155.230 121.370 157.390 ;
        RECT 121.850 155.230 122.200 157.390 ;
        RECT 122.680 155.230 123.030 157.390 ;
        RECT 123.510 155.230 123.860 157.390 ;
        RECT 124.340 155.230 124.690 157.390 ;
        RECT 125.170 155.230 125.520 157.390 ;
        RECT 126.000 155.230 126.350 157.390 ;
        RECT 126.830 155.230 127.180 157.390 ;
        RECT 127.660 155.230 128.010 157.390 ;
        RECT 128.490 155.230 128.840 157.390 ;
        RECT 129.320 155.230 129.670 157.390 ;
        RECT 130.150 155.230 130.500 157.390 ;
        RECT 130.980 155.230 131.330 157.390 ;
        RECT 131.810 155.230 132.160 157.390 ;
        RECT 132.640 155.230 132.990 157.390 ;
        RECT 133.470 155.230 133.820 157.390 ;
        RECT 134.300 155.230 134.650 157.390 ;
        RECT 135.130 155.230 135.480 157.390 ;
        RECT 135.960 155.230 136.310 157.390 ;
        RECT 136.790 155.230 137.140 157.390 ;
        RECT 137.620 155.230 137.970 157.390 ;
        RECT 138.450 155.230 138.800 157.390 ;
        RECT 139.280 155.230 139.630 157.390 ;
        RECT 140.110 155.230 140.460 157.390 ;
        RECT 140.940 155.230 141.290 157.390 ;
        RECT 141.770 155.230 142.120 157.390 ;
        RECT 142.600 155.230 142.950 157.390 ;
        RECT 143.430 155.230 143.780 157.390 ;
        RECT 144.260 155.230 144.610 157.390 ;
        RECT 145.090 155.230 145.440 157.390 ;
        RECT 145.920 155.230 146.270 157.390 ;
        RECT 146.750 155.230 147.100 157.390 ;
        RECT 147.580 155.230 147.930 157.390 ;
        RECT 148.410 155.230 148.760 157.390 ;
        RECT 149.240 155.230 149.590 157.390 ;
        RECT 150.070 155.230 150.420 157.390 ;
        RECT 150.900 155.230 151.250 157.390 ;
        RECT 151.730 155.230 152.080 157.390 ;
        RECT 152.560 155.230 152.910 157.390 ;
        RECT 153.390 155.230 153.740 157.390 ;
        RECT 154.220 155.230 154.570 157.390 ;
        RECT 155.050 155.230 155.400 157.390 ;
        RECT 155.880 155.230 156.230 157.390 ;
        RECT 156.710 155.230 157.060 157.390 ;
        RECT 157.540 155.230 157.890 157.390 ;
        RECT 158.370 155.230 158.720 157.390 ;
        RECT 159.200 155.230 159.550 157.390 ;
        RECT 160.030 155.230 160.380 157.390 ;
        RECT 160.860 155.230 161.210 157.390 ;
        RECT 161.690 155.230 162.040 157.390 ;
        RECT 162.520 155.230 162.870 157.390 ;
        RECT 163.350 155.230 163.700 157.390 ;
        RECT 164.180 155.230 164.530 157.390 ;
        RECT 165.010 155.230 165.360 157.390 ;
        RECT 165.840 155.230 166.190 157.390 ;
        RECT 166.670 155.230 167.020 157.390 ;
        RECT 167.500 155.230 167.850 157.390 ;
        RECT 168.330 155.230 168.680 157.390 ;
        RECT 169.160 155.230 169.510 157.390 ;
        RECT 169.990 155.230 170.340 157.390 ;
        RECT 170.820 155.230 171.170 157.390 ;
        RECT 171.650 155.230 172.000 157.390 ;
        RECT 172.480 155.230 172.830 157.390 ;
        RECT 173.310 155.230 173.660 157.390 ;
        RECT 174.140 155.230 174.490 157.390 ;
        RECT 174.970 155.230 175.320 157.390 ;
        RECT 175.800 155.230 176.150 157.390 ;
        RECT 176.630 155.230 176.980 157.390 ;
        RECT 177.460 155.230 177.810 157.390 ;
        RECT 178.290 155.230 178.640 157.390 ;
        RECT 179.120 155.230 179.470 157.390 ;
        RECT 179.950 155.230 180.300 157.390 ;
        RECT 180.780 155.230 181.130 157.390 ;
        RECT 181.610 155.230 181.960 157.390 ;
        RECT 182.440 155.230 182.790 157.390 ;
        RECT 183.270 155.230 183.620 157.390 ;
        RECT 184.100 155.230 184.450 157.390 ;
        RECT 184.930 155.230 185.280 157.390 ;
        RECT 185.760 155.230 186.110 157.390 ;
        RECT 186.590 155.230 186.940 157.390 ;
        RECT 187.420 155.230 187.770 157.390 ;
        RECT 188.250 155.230 188.600 157.390 ;
        RECT 189.080 155.230 189.430 157.390 ;
        RECT 189.910 155.230 190.260 157.390 ;
        RECT 190.740 155.230 191.090 157.390 ;
        RECT 191.570 155.230 191.920 157.390 ;
        RECT 192.400 155.230 192.750 157.390 ;
        RECT 193.230 155.230 193.580 157.390 ;
        RECT 194.060 155.230 194.410 157.390 ;
        RECT 194.890 155.230 195.240 157.390 ;
        RECT 195.720 155.230 196.070 157.390 ;
        RECT 196.550 155.230 196.900 157.390 ;
        RECT 197.380 155.230 197.730 157.390 ;
        RECT 198.210 155.230 198.560 157.390 ;
        RECT 199.040 155.230 199.390 157.390 ;
        RECT 199.870 155.230 200.220 157.390 ;
        RECT 200.700 155.230 201.050 157.390 ;
        RECT 201.530 155.230 201.880 157.390 ;
        RECT 202.360 155.230 202.710 157.390 ;
        RECT 203.190 155.230 203.540 157.390 ;
        RECT 204.020 155.230 204.370 157.390 ;
        RECT 204.850 155.230 205.200 157.390 ;
        RECT 205.680 155.230 206.030 157.390 ;
        RECT 206.510 155.230 206.860 157.390 ;
        RECT 207.340 155.230 207.690 157.390 ;
        RECT 208.170 155.230 208.520 157.390 ;
        RECT 209.000 155.230 209.350 157.390 ;
        RECT 209.830 155.230 210.180 157.390 ;
        RECT 210.660 155.230 211.010 157.390 ;
        RECT 211.490 155.230 211.840 157.390 ;
        RECT 212.320 154.000 228.050 157.870 ;
        RECT 97.780 151.230 98.130 153.390 ;
        RECT 98.610 151.230 98.960 153.390 ;
        RECT 99.440 151.230 99.790 153.390 ;
        RECT 100.270 151.230 100.620 153.390 ;
        RECT 101.100 151.230 101.450 153.390 ;
        RECT 101.930 151.230 102.280 153.390 ;
        RECT 102.760 151.230 103.110 153.390 ;
        RECT 103.590 151.230 103.940 153.390 ;
        RECT 104.420 151.230 104.770 153.390 ;
        RECT 105.250 151.230 105.600 153.390 ;
        RECT 106.080 151.230 106.430 153.390 ;
        RECT 106.910 151.230 107.260 153.390 ;
        RECT 107.740 151.230 108.090 153.390 ;
        RECT 108.570 151.230 108.920 153.390 ;
        RECT 109.400 151.230 109.750 153.390 ;
        RECT 110.230 151.230 110.580 153.390 ;
        RECT 111.060 151.230 111.410 153.390 ;
        RECT 111.890 151.230 112.240 153.390 ;
        RECT 112.720 151.230 113.070 153.390 ;
        RECT 113.550 151.230 113.900 153.390 ;
        RECT 114.380 151.230 114.730 153.390 ;
        RECT 115.210 151.230 115.560 153.390 ;
        RECT 116.040 151.230 116.390 153.390 ;
        RECT 116.870 151.230 117.220 153.390 ;
        RECT 117.700 151.230 118.050 153.390 ;
        RECT 118.530 151.230 118.880 153.390 ;
        RECT 119.360 151.230 119.710 153.390 ;
        RECT 120.190 151.230 120.540 153.390 ;
        RECT 121.020 151.230 121.370 153.390 ;
        RECT 121.850 151.230 122.200 153.390 ;
        RECT 122.680 151.230 123.030 153.390 ;
        RECT 123.510 151.230 123.860 153.390 ;
        RECT 124.340 151.230 124.690 153.390 ;
        RECT 125.170 151.230 125.520 153.390 ;
        RECT 126.000 151.230 126.350 153.390 ;
        RECT 126.830 151.230 127.180 153.390 ;
        RECT 127.660 151.230 128.010 153.390 ;
        RECT 128.490 151.230 128.840 153.390 ;
        RECT 129.320 151.230 129.670 153.390 ;
        RECT 130.150 151.230 130.500 153.390 ;
        RECT 130.980 151.230 131.330 153.390 ;
        RECT 131.810 151.230 132.160 153.390 ;
        RECT 132.640 151.230 132.990 153.390 ;
        RECT 133.470 151.230 133.820 153.390 ;
        RECT 134.300 151.230 134.650 153.390 ;
        RECT 135.130 151.230 135.480 153.390 ;
        RECT 135.960 151.230 136.310 153.390 ;
        RECT 136.790 151.230 137.140 153.390 ;
        RECT 137.620 151.230 137.970 153.390 ;
        RECT 138.450 151.230 138.800 153.390 ;
        RECT 139.280 151.230 139.630 153.390 ;
        RECT 140.110 151.230 140.460 153.390 ;
        RECT 140.940 151.230 141.290 153.390 ;
        RECT 141.770 151.230 142.120 153.390 ;
        RECT 142.600 151.230 142.950 153.390 ;
        RECT 143.430 151.230 143.780 153.390 ;
        RECT 144.260 151.230 144.610 153.390 ;
        RECT 145.090 151.230 145.440 153.390 ;
        RECT 145.920 151.230 146.270 153.390 ;
        RECT 146.750 151.230 147.100 153.390 ;
        RECT 147.580 151.230 147.930 153.390 ;
        RECT 148.410 151.230 148.760 153.390 ;
        RECT 149.240 151.230 149.590 153.390 ;
        RECT 150.070 151.230 150.420 153.390 ;
        RECT 150.900 151.230 151.250 153.390 ;
        RECT 151.730 151.230 152.080 153.390 ;
        RECT 152.560 151.230 152.910 153.390 ;
        RECT 153.390 151.230 153.740 153.390 ;
        RECT 154.220 151.230 154.570 153.390 ;
        RECT 155.050 151.230 155.400 153.390 ;
        RECT 155.880 151.230 156.230 153.390 ;
        RECT 156.710 151.230 157.060 153.390 ;
        RECT 157.540 151.230 157.890 153.390 ;
        RECT 158.370 151.230 158.720 153.390 ;
        RECT 159.200 151.230 159.550 153.390 ;
        RECT 160.030 151.230 160.380 153.390 ;
        RECT 160.860 151.230 161.210 153.390 ;
        RECT 161.690 151.230 162.040 153.390 ;
        RECT 162.520 151.230 162.870 153.390 ;
        RECT 163.350 151.230 163.700 153.390 ;
        RECT 164.180 151.230 164.530 153.390 ;
        RECT 165.010 151.230 165.360 153.390 ;
        RECT 165.840 151.230 166.190 153.390 ;
        RECT 166.670 151.230 167.020 153.390 ;
        RECT 167.500 151.230 167.850 153.390 ;
        RECT 168.330 151.230 168.680 153.390 ;
        RECT 169.160 151.230 169.510 153.390 ;
        RECT 169.990 151.230 170.340 153.390 ;
        RECT 170.820 151.230 171.170 153.390 ;
        RECT 171.650 151.230 172.000 153.390 ;
        RECT 172.480 151.230 172.830 153.390 ;
        RECT 173.310 151.230 173.660 153.390 ;
        RECT 174.140 151.230 174.490 153.390 ;
        RECT 174.970 151.230 175.320 153.390 ;
        RECT 175.800 151.230 176.150 153.390 ;
        RECT 176.630 151.230 176.980 153.390 ;
        RECT 177.460 151.230 177.810 153.390 ;
        RECT 178.290 151.230 178.640 153.390 ;
        RECT 179.120 151.230 179.470 153.390 ;
        RECT 179.950 151.230 180.300 153.390 ;
        RECT 180.780 151.230 181.130 153.390 ;
        RECT 181.610 151.230 181.960 153.390 ;
        RECT 182.440 151.230 182.790 153.390 ;
        RECT 183.270 151.230 183.620 153.390 ;
        RECT 184.100 151.230 184.450 153.390 ;
        RECT 184.930 151.230 185.280 153.390 ;
        RECT 185.760 151.230 186.110 153.390 ;
        RECT 186.590 151.230 186.940 153.390 ;
        RECT 187.420 151.230 187.770 153.390 ;
        RECT 188.250 151.230 188.600 153.390 ;
        RECT 189.080 151.230 189.430 153.390 ;
        RECT 189.910 151.230 190.260 153.390 ;
        RECT 190.740 151.230 191.090 153.390 ;
        RECT 191.570 151.230 191.920 153.390 ;
        RECT 192.400 151.230 192.750 153.390 ;
        RECT 193.230 151.230 193.580 153.390 ;
        RECT 194.060 151.230 194.410 153.390 ;
        RECT 194.890 151.230 195.240 153.390 ;
        RECT 195.720 151.230 196.070 153.390 ;
        RECT 196.550 151.230 196.900 153.390 ;
        RECT 197.380 151.230 197.730 153.390 ;
        RECT 198.210 151.230 198.560 153.390 ;
        RECT 199.040 151.230 199.390 153.390 ;
        RECT 199.870 151.230 200.220 153.390 ;
        RECT 200.700 151.230 201.050 153.390 ;
        RECT 201.530 151.230 201.880 153.390 ;
        RECT 202.360 151.230 202.710 153.390 ;
        RECT 203.190 151.230 203.540 153.390 ;
        RECT 204.020 151.230 204.370 153.390 ;
        RECT 204.850 151.230 205.200 153.390 ;
        RECT 205.680 151.230 206.030 153.390 ;
        RECT 206.510 151.230 206.860 153.390 ;
        RECT 207.340 151.230 207.690 153.390 ;
        RECT 208.170 151.230 208.520 153.390 ;
        RECT 209.000 151.230 209.350 153.390 ;
        RECT 209.830 151.230 210.180 153.390 ;
        RECT 210.660 151.230 211.010 153.390 ;
        RECT 211.490 151.230 211.840 153.390 ;
        RECT 212.320 150.750 212.675 154.000 ;
        RECT 75.275 150.600 212.675 150.750 ;
        RECT 215.625 153.550 228.050 154.000 ;
        RECT 231.045 158.645 271.250 158.995 ;
        RECT 231.045 158.640 249.805 158.645 ;
        RECT 231.045 157.900 231.400 158.640 ;
        RECT 231.670 158.120 232.195 158.445 ;
        RECT 233.495 158.120 234.020 158.445 ;
        RECT 231.800 157.900 231.970 157.915 ;
        RECT 232.280 157.900 232.450 157.915 ;
        RECT 231.045 154.875 232.475 157.900 ;
        RECT 232.760 154.875 232.930 157.915 ;
        RECT 233.240 157.900 233.410 157.915 ;
        RECT 233.720 157.900 233.890 157.915 ;
        RECT 234.290 157.900 236.000 158.640 ;
        RECT 236.270 158.120 236.795 158.445 ;
        RECT 238.095 158.120 238.620 158.445 ;
        RECT 236.400 157.900 236.570 157.915 ;
        RECT 236.880 157.900 237.050 157.915 ;
        RECT 233.225 154.875 237.075 157.900 ;
        RECT 237.360 154.875 237.530 157.915 ;
        RECT 237.840 157.900 238.010 157.915 ;
        RECT 238.320 157.900 238.490 157.915 ;
        RECT 238.890 157.900 240.600 158.640 ;
        RECT 242.570 158.120 242.945 158.445 ;
        RECT 241.000 157.900 241.170 157.915 ;
        RECT 241.480 157.900 241.650 157.915 ;
        RECT 237.825 154.875 241.675 157.900 ;
        RECT 241.960 154.875 242.130 157.915 ;
        RECT 242.440 157.900 242.610 157.915 ;
        RECT 242.920 157.900 243.090 157.915 ;
        RECT 243.490 157.900 245.200 158.640 ;
        RECT 245.470 158.120 245.995 158.445 ;
        RECT 247.295 158.120 247.820 158.445 ;
        RECT 248.090 157.925 249.805 158.640 ;
        RECT 250.080 158.125 250.580 158.450 ;
        RECT 253.830 158.125 254.330 158.450 ;
        RECT 254.605 157.925 271.250 158.645 ;
        RECT 245.600 157.900 245.770 157.915 ;
        RECT 246.080 157.900 246.250 157.915 ;
        RECT 242.425 154.875 246.275 157.900 ;
        RECT 246.560 154.875 246.730 157.915 ;
        RECT 247.040 157.900 247.210 157.915 ;
        RECT 247.520 157.900 247.690 157.915 ;
        RECT 248.090 157.900 250.875 157.925 ;
        RECT 247.025 154.875 250.875 157.900 ;
        RECT 251.160 154.880 251.330 157.920 ;
        RECT 251.640 154.880 251.810 157.920 ;
        RECT 252.120 154.880 252.290 157.920 ;
        RECT 252.600 154.880 252.770 157.920 ;
        RECT 253.080 154.880 253.250 157.920 ;
        RECT 253.525 154.875 271.250 157.925 ;
        RECT 231.045 154.150 231.400 154.875 ;
        RECT 232.445 154.320 233.245 154.695 ;
        RECT 234.290 154.150 236.000 154.875 ;
        RECT 237.045 154.320 237.845 154.695 ;
        RECT 238.890 154.150 240.600 154.875 ;
        RECT 242.095 154.320 242.470 154.695 ;
        RECT 243.490 154.150 245.200 154.875 ;
        RECT 246.245 154.320 247.045 154.695 ;
        RECT 248.090 154.155 249.805 154.875 ;
        RECT 250.830 154.325 253.580 154.700 ;
        RECT 254.605 154.155 271.250 154.875 ;
        RECT 248.090 154.150 271.250 154.155 ;
        RECT 231.045 153.800 271.250 154.150 ;
        RECT 231.045 153.795 234.645 153.800 ;
        RECT 235.645 153.795 239.245 153.800 ;
        RECT 240.245 153.795 243.845 153.800 ;
        RECT 244.845 153.795 248.445 153.800 ;
        RECT 215.625 153.200 254.955 153.550 ;
        RECT 215.625 152.525 231.405 153.200 ;
        RECT 232.450 152.700 233.250 153.025 ;
        RECT 234.295 152.525 236.005 153.200 ;
        RECT 237.050 152.700 237.850 153.025 ;
        RECT 238.895 152.525 240.605 153.200 ;
        RECT 242.100 152.700 242.475 153.025 ;
        RECT 243.495 152.525 245.205 153.200 ;
        RECT 246.250 152.700 247.050 153.025 ;
        RECT 248.095 152.525 249.805 153.200 ;
        RECT 250.830 152.700 253.580 153.025 ;
        RECT 254.605 152.525 254.955 153.200 ;
        RECT 215.625 151.475 232.475 152.525 ;
        RECT 232.765 151.480 232.935 152.520 ;
        RECT 233.225 151.475 237.075 152.525 ;
        RECT 237.365 151.480 237.535 152.520 ;
        RECT 237.825 151.475 241.675 152.525 ;
        RECT 241.965 151.480 242.135 152.520 ;
        RECT 242.425 151.475 246.275 152.525 ;
        RECT 246.565 151.480 246.735 152.520 ;
        RECT 247.025 151.475 250.875 152.525 ;
        RECT 251.160 151.480 251.330 152.520 ;
        RECT 251.640 151.480 251.810 152.520 ;
        RECT 252.120 151.480 252.290 152.520 ;
        RECT 252.600 151.480 252.770 152.520 ;
        RECT 253.080 151.480 253.250 152.520 ;
        RECT 253.525 151.475 254.955 152.525 ;
        RECT 215.625 150.800 231.405 151.475 ;
        RECT 231.675 150.975 232.200 151.300 ;
        RECT 233.500 150.975 234.025 151.300 ;
        RECT 234.295 150.800 236.005 151.475 ;
        RECT 236.275 150.975 236.800 151.300 ;
        RECT 238.100 150.975 238.625 151.300 ;
        RECT 238.895 150.800 240.605 151.475 ;
        RECT 242.575 150.975 242.950 151.300 ;
        RECT 243.495 150.800 245.205 151.475 ;
        RECT 245.475 150.975 246.000 151.300 ;
        RECT 247.300 150.975 247.825 151.300 ;
        RECT 248.095 150.800 249.805 151.475 ;
        RECT 250.080 150.975 250.580 151.300 ;
        RECT 253.830 150.975 254.330 151.300 ;
        RECT 254.605 150.800 254.955 151.475 ;
        RECT 215.625 150.600 254.955 150.800 ;
        RECT 75.275 150.580 212.490 150.600 ;
        RECT 75.275 150.575 97.300 150.580 ;
        RECT 226.800 150.450 254.955 150.600 ;
        RECT 256.625 152.940 271.250 153.800 ;
        RECT 65.075 148.250 70.925 149.825 ;
        RECT 75.280 147.560 226.130 149.895 ;
        RECT 75.280 146.835 76.030 147.560 ;
        RECT 76.260 147.050 77.260 147.220 ;
        RECT 82.710 147.050 83.710 147.220 ;
        RECT 83.930 146.835 86.805 147.560 ;
        RECT 87.010 147.050 88.010 147.220 ;
        RECT 96.040 147.050 97.040 147.220 ;
        RECT 97.255 146.835 100.130 147.560 ;
        RECT 100.335 147.050 101.335 147.220 ;
        RECT 109.365 147.050 110.365 147.220 ;
        RECT 110.580 146.835 113.430 147.560 ;
        RECT 113.660 147.050 114.660 147.220 ;
        RECT 120.110 147.050 121.110 147.220 ;
        RECT 121.330 146.835 124.205 147.560 ;
        RECT 124.410 147.050 125.410 147.220 ;
        RECT 133.440 147.050 134.440 147.220 ;
        RECT 134.655 146.835 137.530 147.560 ;
        RECT 137.735 147.050 138.735 147.220 ;
        RECT 146.765 147.050 147.765 147.220 ;
        RECT 147.980 146.835 150.855 147.560 ;
        RECT 151.060 147.050 152.060 147.220 ;
        RECT 160.090 147.050 161.090 147.220 ;
        RECT 161.305 146.835 164.180 147.560 ;
        RECT 164.385 147.050 165.385 147.220 ;
        RECT 173.415 147.050 174.415 147.220 ;
        RECT 174.630 146.835 177.505 147.560 ;
        RECT 177.710 147.050 178.710 147.220 ;
        RECT 186.740 147.050 187.740 147.220 ;
        RECT 187.955 146.835 190.805 147.560 ;
        RECT 191.035 147.050 192.035 147.220 ;
        RECT 197.485 147.050 198.485 147.220 ;
        RECT 198.705 146.835 201.580 147.560 ;
        RECT 201.785 147.050 202.785 147.220 ;
        RECT 210.815 147.050 211.815 147.220 ;
        RECT 212.030 146.835 214.905 147.560 ;
        RECT 215.110 147.050 216.110 147.220 ;
        RECT 224.140 147.050 225.140 147.220 ;
        RECT 225.355 146.835 226.130 147.560 ;
        RECT 75.280 137.795 76.200 146.835 ;
        RECT 77.320 137.795 77.490 146.835 ;
        RECT 78.610 137.795 78.780 146.835 ;
        RECT 79.900 137.795 80.070 146.835 ;
        RECT 81.190 137.795 81.360 146.835 ;
        RECT 82.480 137.795 82.650 146.835 ;
        RECT 83.770 137.795 86.950 146.835 ;
        RECT 88.070 137.795 88.240 146.835 ;
        RECT 89.360 137.795 89.530 146.835 ;
        RECT 90.650 137.795 90.820 146.835 ;
        RECT 91.940 137.795 92.110 146.835 ;
        RECT 93.230 137.795 93.400 146.835 ;
        RECT 94.520 137.795 94.690 146.835 ;
        RECT 95.810 137.795 95.980 146.835 ;
        RECT 97.100 137.795 100.275 146.835 ;
        RECT 101.395 137.795 101.565 146.835 ;
        RECT 102.685 137.795 102.855 146.835 ;
        RECT 103.975 137.795 104.145 146.835 ;
        RECT 105.265 137.795 105.435 146.835 ;
        RECT 106.555 137.795 106.725 146.835 ;
        RECT 107.845 137.795 108.015 146.835 ;
        RECT 109.135 137.795 109.305 146.835 ;
        RECT 110.425 137.795 113.600 146.835 ;
        RECT 114.720 137.795 114.890 146.835 ;
        RECT 116.010 137.795 116.180 146.835 ;
        RECT 117.300 137.795 117.470 146.835 ;
        RECT 118.590 137.795 118.760 146.835 ;
        RECT 119.880 137.795 120.050 146.835 ;
        RECT 121.170 137.795 124.350 146.835 ;
        RECT 125.470 137.795 125.640 146.835 ;
        RECT 126.760 137.795 126.930 146.835 ;
        RECT 128.050 137.795 128.220 146.835 ;
        RECT 129.340 137.795 129.510 146.835 ;
        RECT 130.630 137.795 130.800 146.835 ;
        RECT 131.920 137.795 132.090 146.835 ;
        RECT 133.210 137.795 133.380 146.835 ;
        RECT 134.500 137.795 137.675 146.835 ;
        RECT 138.795 137.795 138.965 146.835 ;
        RECT 140.085 137.795 140.255 146.835 ;
        RECT 141.375 137.795 141.545 146.835 ;
        RECT 142.665 137.795 142.835 146.835 ;
        RECT 143.955 137.795 144.125 146.835 ;
        RECT 145.245 137.795 145.415 146.835 ;
        RECT 146.535 137.795 146.705 146.835 ;
        RECT 147.825 137.795 151.000 146.835 ;
        RECT 152.120 137.795 152.290 146.835 ;
        RECT 153.410 137.795 153.580 146.835 ;
        RECT 154.700 137.795 154.870 146.835 ;
        RECT 155.990 137.795 156.160 146.835 ;
        RECT 157.280 137.795 157.450 146.835 ;
        RECT 158.570 137.795 158.740 146.835 ;
        RECT 159.860 137.795 160.030 146.835 ;
        RECT 161.150 137.795 164.325 146.835 ;
        RECT 165.445 137.795 165.615 146.835 ;
        RECT 166.735 137.795 166.905 146.835 ;
        RECT 168.025 137.795 168.195 146.835 ;
        RECT 169.315 137.795 169.485 146.835 ;
        RECT 170.605 137.795 170.775 146.835 ;
        RECT 171.895 137.795 172.065 146.835 ;
        RECT 173.185 137.795 173.355 146.835 ;
        RECT 174.475 137.795 177.650 146.835 ;
        RECT 178.770 137.795 178.940 146.835 ;
        RECT 180.060 137.795 180.230 146.835 ;
        RECT 181.350 137.795 181.520 146.835 ;
        RECT 182.640 137.795 182.810 146.835 ;
        RECT 183.930 137.795 184.100 146.835 ;
        RECT 185.220 137.795 185.390 146.835 ;
        RECT 186.510 137.795 186.680 146.835 ;
        RECT 187.800 137.795 190.975 146.835 ;
        RECT 192.095 137.795 192.265 146.835 ;
        RECT 193.385 137.795 193.555 146.835 ;
        RECT 194.675 137.795 194.845 146.835 ;
        RECT 195.965 137.795 196.135 146.835 ;
        RECT 197.255 137.795 197.425 146.835 ;
        RECT 198.545 137.795 201.725 146.835 ;
        RECT 202.845 137.795 203.015 146.835 ;
        RECT 204.135 137.795 204.305 146.835 ;
        RECT 205.425 137.795 205.595 146.835 ;
        RECT 206.715 137.795 206.885 146.835 ;
        RECT 208.005 137.795 208.175 146.835 ;
        RECT 209.295 137.795 209.465 146.835 ;
        RECT 210.585 137.795 210.755 146.835 ;
        RECT 211.875 137.795 215.050 146.835 ;
        RECT 216.170 137.795 216.340 146.835 ;
        RECT 217.460 137.795 217.630 146.835 ;
        RECT 218.750 137.795 218.920 146.835 ;
        RECT 220.040 137.795 220.210 146.835 ;
        RECT 221.330 137.795 221.500 146.835 ;
        RECT 222.620 137.795 222.790 146.835 ;
        RECT 223.910 137.795 224.080 146.835 ;
        RECT 225.200 137.795 226.130 146.835 ;
        RECT 75.280 137.195 76.030 137.795 ;
        RECT 77.550 137.410 78.550 137.580 ;
        RECT 78.840 137.410 79.840 137.580 ;
        RECT 80.130 137.410 81.130 137.580 ;
        RECT 81.420 137.410 82.420 137.580 ;
        RECT 83.930 137.195 86.805 137.795 ;
        RECT 88.300 137.410 89.300 137.580 ;
        RECT 89.590 137.410 90.590 137.580 ;
        RECT 90.880 137.410 91.880 137.580 ;
        RECT 92.170 137.410 93.170 137.580 ;
        RECT 93.460 137.410 94.460 137.580 ;
        RECT 94.750 137.410 95.750 137.580 ;
        RECT 97.255 137.195 100.130 137.795 ;
        RECT 101.625 137.410 102.625 137.580 ;
        RECT 102.915 137.410 103.915 137.580 ;
        RECT 104.205 137.410 105.205 137.580 ;
        RECT 105.495 137.410 106.495 137.580 ;
        RECT 106.785 137.410 107.785 137.580 ;
        RECT 108.075 137.410 109.075 137.580 ;
        RECT 110.580 137.195 113.430 137.795 ;
        RECT 114.950 137.410 115.950 137.580 ;
        RECT 116.240 137.410 117.240 137.580 ;
        RECT 117.530 137.410 118.530 137.580 ;
        RECT 118.820 137.410 119.820 137.580 ;
        RECT 121.330 137.195 124.205 137.795 ;
        RECT 125.700 137.410 126.700 137.580 ;
        RECT 126.990 137.410 127.990 137.580 ;
        RECT 128.280 137.410 129.280 137.580 ;
        RECT 129.570 137.410 130.570 137.580 ;
        RECT 130.860 137.410 131.860 137.580 ;
        RECT 132.150 137.410 133.150 137.580 ;
        RECT 134.655 137.195 137.530 137.795 ;
        RECT 139.025 137.410 140.025 137.580 ;
        RECT 140.315 137.410 141.315 137.580 ;
        RECT 141.605 137.410 142.605 137.580 ;
        RECT 142.895 137.410 143.895 137.580 ;
        RECT 144.185 137.410 145.185 137.580 ;
        RECT 145.475 137.410 146.475 137.580 ;
        RECT 147.980 137.195 150.855 137.795 ;
        RECT 152.350 137.410 153.350 137.580 ;
        RECT 153.640 137.410 154.640 137.580 ;
        RECT 154.930 137.410 155.930 137.580 ;
        RECT 156.220 137.410 157.220 137.580 ;
        RECT 157.510 137.410 158.510 137.580 ;
        RECT 158.800 137.410 159.800 137.580 ;
        RECT 161.305 137.195 164.180 137.795 ;
        RECT 165.675 137.410 166.675 137.580 ;
        RECT 166.965 137.410 167.965 137.580 ;
        RECT 168.255 137.410 169.255 137.580 ;
        RECT 169.545 137.410 170.545 137.580 ;
        RECT 170.835 137.410 171.835 137.580 ;
        RECT 172.125 137.410 173.125 137.580 ;
        RECT 174.630 137.195 177.505 137.795 ;
        RECT 179.000 137.410 180.000 137.580 ;
        RECT 180.290 137.410 181.290 137.580 ;
        RECT 181.580 137.410 182.580 137.580 ;
        RECT 182.870 137.410 183.870 137.580 ;
        RECT 184.160 137.410 185.160 137.580 ;
        RECT 185.450 137.410 186.450 137.580 ;
        RECT 187.955 137.195 190.805 137.795 ;
        RECT 192.325 137.410 193.325 137.580 ;
        RECT 193.615 137.410 194.615 137.580 ;
        RECT 194.905 137.410 195.905 137.580 ;
        RECT 196.195 137.410 197.195 137.580 ;
        RECT 198.705 137.195 201.580 137.795 ;
        RECT 203.075 137.410 204.075 137.580 ;
        RECT 204.365 137.410 205.365 137.580 ;
        RECT 205.655 137.410 206.655 137.580 ;
        RECT 206.945 137.410 207.945 137.580 ;
        RECT 208.235 137.410 209.235 137.580 ;
        RECT 209.525 137.410 210.525 137.580 ;
        RECT 212.030 137.195 214.905 137.795 ;
        RECT 216.400 137.410 217.400 137.580 ;
        RECT 217.690 137.410 218.690 137.580 ;
        RECT 218.980 137.410 219.980 137.580 ;
        RECT 220.270 137.410 221.270 137.580 ;
        RECT 221.560 137.410 222.560 137.580 ;
        RECT 222.850 137.410 223.850 137.580 ;
        RECT 225.355 137.195 226.130 137.795 ;
        RECT 72.725 136.075 73.450 137.175 ;
        RECT 75.280 136.900 226.130 137.195 ;
        RECT 75.280 136.895 76.030 136.900 ;
        RECT 83.930 136.895 86.805 136.900 ;
        RECT 97.255 136.895 100.130 136.900 ;
        RECT 110.580 136.895 113.430 136.900 ;
        RECT 121.330 136.895 124.205 136.900 ;
        RECT 134.655 136.895 137.530 136.900 ;
        RECT 147.980 136.895 150.855 136.900 ;
        RECT 161.305 136.895 164.180 136.900 ;
        RECT 174.630 136.895 177.505 136.900 ;
        RECT 187.955 136.895 190.805 136.900 ;
        RECT 198.705 136.895 201.580 136.900 ;
        RECT 212.030 136.895 214.905 136.900 ;
        RECT 225.355 136.895 226.130 136.900 ;
        RECT 226.800 144.250 228.050 150.450 ;
        RECT 231.050 149.700 233.700 149.705 ;
        RECT 231.050 149.350 254.955 149.700 ;
        RECT 231.050 144.860 231.425 149.350 ;
        RECT 233.325 149.345 254.955 149.350 ;
        RECT 233.325 149.340 249.805 149.345 ;
        RECT 231.950 148.805 232.800 149.180 ;
        RECT 231.810 145.585 231.980 148.625 ;
        RECT 232.290 145.585 232.460 148.625 ;
        RECT 232.770 145.585 232.940 148.625 ;
        RECT 233.325 148.600 236.000 149.340 ;
        RECT 236.270 148.820 236.795 149.145 ;
        RECT 238.095 148.820 238.620 149.145 ;
        RECT 236.400 148.600 236.570 148.615 ;
        RECT 236.880 148.600 237.050 148.615 ;
        RECT 233.325 145.575 237.075 148.600 ;
        RECT 237.360 145.575 237.530 148.615 ;
        RECT 237.840 148.600 238.010 148.615 ;
        RECT 238.320 148.600 238.490 148.615 ;
        RECT 238.890 148.600 240.600 149.340 ;
        RECT 242.570 148.820 242.945 149.145 ;
        RECT 241.000 148.600 241.170 148.615 ;
        RECT 241.480 148.600 241.650 148.615 ;
        RECT 237.825 145.575 241.675 148.600 ;
        RECT 241.960 145.575 242.130 148.615 ;
        RECT 242.440 148.600 242.610 148.615 ;
        RECT 242.920 148.600 243.090 148.615 ;
        RECT 243.490 148.600 245.200 149.340 ;
        RECT 245.470 148.820 245.995 149.145 ;
        RECT 247.295 148.820 247.820 149.145 ;
        RECT 248.090 148.625 249.805 149.340 ;
        RECT 250.080 148.825 250.580 149.150 ;
        RECT 253.830 148.825 254.330 149.150 ;
        RECT 254.605 148.625 254.955 149.345 ;
        RECT 245.600 148.600 245.770 148.615 ;
        RECT 246.080 148.600 246.250 148.615 ;
        RECT 242.425 145.575 246.275 148.600 ;
        RECT 246.560 145.575 246.730 148.615 ;
        RECT 247.040 148.600 247.210 148.615 ;
        RECT 247.520 148.600 247.690 148.615 ;
        RECT 248.090 148.600 250.875 148.625 ;
        RECT 247.025 145.575 250.875 148.600 ;
        RECT 251.160 145.580 251.330 148.620 ;
        RECT 251.640 145.580 251.810 148.620 ;
        RECT 252.120 145.580 252.290 148.620 ;
        RECT 252.600 145.580 252.770 148.620 ;
        RECT 253.080 145.580 253.250 148.620 ;
        RECT 253.525 145.575 254.955 148.625 ;
        RECT 256.625 148.450 256.975 152.940 ;
        RECT 257.540 152.395 259.290 152.770 ;
        RECT 268.590 152.395 270.340 152.770 ;
        RECT 257.375 149.175 257.545 152.215 ;
        RECT 257.855 149.175 258.025 152.215 ;
        RECT 258.335 149.175 258.505 152.215 ;
        RECT 258.815 149.175 258.985 152.215 ;
        RECT 259.295 149.175 259.465 152.215 ;
        RECT 259.775 149.175 259.945 152.215 ;
        RECT 260.255 149.175 260.425 152.215 ;
        RECT 260.735 149.175 260.905 152.215 ;
        RECT 261.215 149.175 261.385 152.215 ;
        RECT 261.695 149.175 261.865 152.215 ;
        RECT 262.175 149.175 262.345 152.215 ;
        RECT 262.655 149.175 262.825 152.215 ;
        RECT 263.135 149.175 263.305 152.215 ;
        RECT 263.615 149.175 263.785 152.215 ;
        RECT 264.095 149.175 264.265 152.215 ;
        RECT 264.575 149.175 264.745 152.215 ;
        RECT 265.055 149.175 265.225 152.215 ;
        RECT 265.535 149.175 265.705 152.215 ;
        RECT 266.015 149.175 266.185 152.215 ;
        RECT 266.495 149.175 266.665 152.215 ;
        RECT 266.975 149.175 267.145 152.215 ;
        RECT 267.455 149.175 267.625 152.215 ;
        RECT 267.935 149.175 268.105 152.215 ;
        RECT 268.415 149.175 268.585 152.215 ;
        RECT 268.895 149.175 269.065 152.215 ;
        RECT 269.375 149.175 269.545 152.215 ;
        RECT 269.855 149.175 270.025 152.215 ;
        RECT 270.335 149.175 270.505 152.215 ;
        RECT 259.465 148.620 268.415 148.995 ;
        RECT 270.900 148.450 271.250 152.940 ;
        RECT 256.625 148.100 271.250 148.450 ;
        RECT 233.325 144.860 236.000 145.575 ;
        RECT 237.045 145.020 237.845 145.395 ;
        RECT 231.050 144.850 236.000 144.860 ;
        RECT 238.890 144.850 240.600 145.575 ;
        RECT 242.095 145.020 242.470 145.395 ;
        RECT 243.490 144.850 245.200 145.575 ;
        RECT 246.245 145.020 247.045 145.395 ;
        RECT 248.090 144.855 249.805 145.575 ;
        RECT 250.830 145.025 253.580 145.400 ;
        RECT 254.605 144.855 254.955 145.575 ;
        RECT 248.090 144.850 254.955 144.855 ;
        RECT 231.050 144.505 254.955 144.850 ;
        RECT 233.325 144.500 254.955 144.505 ;
        RECT 256.625 147.500 271.250 147.850 ;
        RECT 256.625 145.100 256.975 147.500 ;
        RECT 257.540 147.000 259.290 147.325 ;
        RECT 268.590 147.000 270.340 147.325 ;
        RECT 257.375 145.780 257.545 146.820 ;
        RECT 257.855 145.780 258.025 146.820 ;
        RECT 258.335 145.780 258.505 146.820 ;
        RECT 258.815 145.780 258.985 146.820 ;
        RECT 259.295 145.780 259.465 146.820 ;
        RECT 259.775 145.780 259.945 146.820 ;
        RECT 260.255 145.780 260.425 146.820 ;
        RECT 260.735 145.780 260.905 146.820 ;
        RECT 261.215 145.780 261.385 146.820 ;
        RECT 261.695 145.780 261.865 146.820 ;
        RECT 262.175 145.780 262.345 146.820 ;
        RECT 262.655 145.780 262.825 146.820 ;
        RECT 263.135 145.780 263.305 146.820 ;
        RECT 263.615 145.780 263.785 146.820 ;
        RECT 264.095 145.780 264.265 146.820 ;
        RECT 264.575 145.780 264.745 146.820 ;
        RECT 265.055 145.780 265.225 146.820 ;
        RECT 265.535 145.780 265.705 146.820 ;
        RECT 266.015 145.780 266.185 146.820 ;
        RECT 266.495 145.780 266.665 146.820 ;
        RECT 266.975 145.780 267.145 146.820 ;
        RECT 267.455 145.780 267.625 146.820 ;
        RECT 267.935 145.780 268.105 146.820 ;
        RECT 268.415 145.780 268.585 146.820 ;
        RECT 268.895 145.780 269.065 146.820 ;
        RECT 269.375 145.780 269.545 146.820 ;
        RECT 269.855 145.780 270.025 146.820 ;
        RECT 270.335 145.780 270.505 146.820 ;
        RECT 259.465 145.275 268.415 145.600 ;
        RECT 270.900 145.100 271.250 147.500 ;
        RECT 235.645 144.495 239.245 144.500 ;
        RECT 240.245 144.495 243.845 144.500 ;
        RECT 244.845 144.495 248.445 144.500 ;
        RECT 256.625 144.250 271.250 145.100 ;
        RECT 226.800 143.900 271.250 144.250 ;
        RECT 226.800 141.500 231.425 143.900 ;
        RECT 233.325 143.225 236.005 143.900 ;
        RECT 237.050 143.400 237.850 143.725 ;
        RECT 238.895 143.225 240.605 143.900 ;
        RECT 242.100 143.400 242.475 143.725 ;
        RECT 243.495 143.225 245.205 143.900 ;
        RECT 246.250 143.400 247.050 143.725 ;
        RECT 248.095 143.225 249.805 143.900 ;
        RECT 250.830 143.400 253.580 143.725 ;
        RECT 254.605 143.225 271.250 143.900 ;
        RECT 231.810 142.180 231.980 143.220 ;
        RECT 232.290 142.180 232.460 143.220 ;
        RECT 232.770 142.180 232.940 143.220 ;
        RECT 233.325 142.175 237.075 143.225 ;
        RECT 237.365 142.180 237.535 143.220 ;
        RECT 237.825 142.175 241.675 143.225 ;
        RECT 241.965 142.180 242.135 143.220 ;
        RECT 242.425 142.175 246.275 143.225 ;
        RECT 246.565 142.180 246.735 143.220 ;
        RECT 247.025 142.175 250.875 143.225 ;
        RECT 251.160 142.180 251.330 143.220 ;
        RECT 251.640 142.180 251.810 143.220 ;
        RECT 252.120 142.180 252.290 143.220 ;
        RECT 252.600 142.180 252.770 143.220 ;
        RECT 253.080 142.180 253.250 143.220 ;
        RECT 253.525 142.175 271.250 143.225 ;
        RECT 231.950 141.675 232.800 142.000 ;
        RECT 233.325 141.500 236.005 142.175 ;
        RECT 236.275 141.675 236.800 142.000 ;
        RECT 238.100 141.675 238.625 142.000 ;
        RECT 238.895 141.500 240.605 142.175 ;
        RECT 242.575 141.675 242.950 142.000 ;
        RECT 243.495 141.500 245.205 142.175 ;
        RECT 245.475 141.675 246.000 142.000 ;
        RECT 247.300 141.675 247.825 142.000 ;
        RECT 248.095 141.500 249.805 142.175 ;
        RECT 250.080 141.675 250.580 142.000 ;
        RECT 253.830 141.675 254.330 142.000 ;
        RECT 254.605 141.500 271.250 142.175 ;
        RECT 226.800 140.300 271.250 141.500 ;
        RECT 75.280 136.045 226.130 136.345 ;
        RECT 75.280 135.490 76.030 136.045 ;
        RECT 77.550 135.660 78.550 135.830 ;
        RECT 78.840 135.660 79.840 135.830 ;
        RECT 80.130 135.660 81.130 135.830 ;
        RECT 81.420 135.660 82.420 135.830 ;
        RECT 83.930 135.490 86.805 136.045 ;
        RECT 88.300 135.660 89.300 135.830 ;
        RECT 89.590 135.660 90.590 135.830 ;
        RECT 90.880 135.660 91.880 135.830 ;
        RECT 92.170 135.660 93.170 135.830 ;
        RECT 93.460 135.660 94.460 135.830 ;
        RECT 94.750 135.660 95.750 135.830 ;
        RECT 97.255 135.490 100.130 136.045 ;
        RECT 101.625 135.660 102.625 135.830 ;
        RECT 102.915 135.660 103.915 135.830 ;
        RECT 104.205 135.660 105.205 135.830 ;
        RECT 105.495 135.660 106.495 135.830 ;
        RECT 106.785 135.660 107.785 135.830 ;
        RECT 108.075 135.660 109.075 135.830 ;
        RECT 110.580 135.490 113.430 136.045 ;
        RECT 114.950 135.660 115.950 135.830 ;
        RECT 116.240 135.660 117.240 135.830 ;
        RECT 117.530 135.660 118.530 135.830 ;
        RECT 118.820 135.660 119.820 135.830 ;
        RECT 121.330 135.490 124.205 136.045 ;
        RECT 125.700 135.660 126.700 135.830 ;
        RECT 126.990 135.660 127.990 135.830 ;
        RECT 128.280 135.660 129.280 135.830 ;
        RECT 129.570 135.660 130.570 135.830 ;
        RECT 130.860 135.660 131.860 135.830 ;
        RECT 132.150 135.660 133.150 135.830 ;
        RECT 134.655 135.490 137.530 136.045 ;
        RECT 139.025 135.660 140.025 135.830 ;
        RECT 140.315 135.660 141.315 135.830 ;
        RECT 141.605 135.660 142.605 135.830 ;
        RECT 142.895 135.660 143.895 135.830 ;
        RECT 144.185 135.660 145.185 135.830 ;
        RECT 145.475 135.660 146.475 135.830 ;
        RECT 147.980 135.490 150.855 136.045 ;
        RECT 152.350 135.660 153.350 135.830 ;
        RECT 153.640 135.660 154.640 135.830 ;
        RECT 154.930 135.660 155.930 135.830 ;
        RECT 156.220 135.660 157.220 135.830 ;
        RECT 157.510 135.660 158.510 135.830 ;
        RECT 158.800 135.660 159.800 135.830 ;
        RECT 161.305 135.490 164.180 136.045 ;
        RECT 165.675 135.660 166.675 135.830 ;
        RECT 166.965 135.660 167.965 135.830 ;
        RECT 168.255 135.660 169.255 135.830 ;
        RECT 169.545 135.660 170.545 135.830 ;
        RECT 170.835 135.660 171.835 135.830 ;
        RECT 172.125 135.660 173.125 135.830 ;
        RECT 174.630 135.490 177.505 136.045 ;
        RECT 179.000 135.660 180.000 135.830 ;
        RECT 180.290 135.660 181.290 135.830 ;
        RECT 181.580 135.660 182.580 135.830 ;
        RECT 182.870 135.660 183.870 135.830 ;
        RECT 184.160 135.660 185.160 135.830 ;
        RECT 185.450 135.660 186.450 135.830 ;
        RECT 187.955 135.490 190.805 136.045 ;
        RECT 192.325 135.660 193.325 135.830 ;
        RECT 193.615 135.660 194.615 135.830 ;
        RECT 194.905 135.660 195.905 135.830 ;
        RECT 196.195 135.660 197.195 135.830 ;
        RECT 198.705 135.490 201.580 136.045 ;
        RECT 203.075 135.660 204.075 135.830 ;
        RECT 204.365 135.660 205.365 135.830 ;
        RECT 205.655 135.660 206.655 135.830 ;
        RECT 206.945 135.660 207.945 135.830 ;
        RECT 208.235 135.660 209.235 135.830 ;
        RECT 209.525 135.660 210.525 135.830 ;
        RECT 212.030 135.490 214.905 136.045 ;
        RECT 216.400 135.660 217.400 135.830 ;
        RECT 217.690 135.660 218.690 135.830 ;
        RECT 218.980 135.660 219.980 135.830 ;
        RECT 220.270 135.660 221.270 135.830 ;
        RECT 221.560 135.660 222.560 135.830 ;
        RECT 222.850 135.660 223.850 135.830 ;
        RECT 225.355 135.500 226.130 136.045 ;
        RECT 226.800 135.500 228.050 140.300 ;
        RECT 231.050 138.145 271.250 139.000 ;
        RECT 225.355 135.490 228.050 135.500 ;
        RECT 75.280 132.450 76.200 135.490 ;
        RECT 77.320 132.450 77.490 135.490 ;
        RECT 78.610 132.450 78.780 135.490 ;
        RECT 79.900 132.450 80.070 135.490 ;
        RECT 81.190 132.450 81.360 135.490 ;
        RECT 82.480 132.450 82.650 135.490 ;
        RECT 83.770 132.450 86.950 135.490 ;
        RECT 88.070 132.450 88.240 135.490 ;
        RECT 89.360 132.450 89.530 135.490 ;
        RECT 90.650 132.450 90.820 135.490 ;
        RECT 91.940 132.450 92.110 135.490 ;
        RECT 93.230 132.450 93.400 135.490 ;
        RECT 94.520 132.450 94.690 135.490 ;
        RECT 95.810 132.450 95.980 135.490 ;
        RECT 97.100 132.450 100.275 135.490 ;
        RECT 101.395 132.450 101.565 135.490 ;
        RECT 102.685 132.450 102.855 135.490 ;
        RECT 103.975 132.450 104.145 135.490 ;
        RECT 105.265 132.450 105.435 135.490 ;
        RECT 106.555 132.450 106.725 135.490 ;
        RECT 107.845 132.450 108.015 135.490 ;
        RECT 109.135 132.450 109.305 135.490 ;
        RECT 110.425 132.450 113.600 135.490 ;
        RECT 114.720 132.450 114.890 135.490 ;
        RECT 116.010 132.450 116.180 135.490 ;
        RECT 117.300 132.450 117.470 135.490 ;
        RECT 118.590 132.450 118.760 135.490 ;
        RECT 119.880 132.450 120.050 135.490 ;
        RECT 121.170 132.450 124.350 135.490 ;
        RECT 125.470 132.450 125.640 135.490 ;
        RECT 126.760 132.450 126.930 135.490 ;
        RECT 128.050 132.450 128.220 135.490 ;
        RECT 129.340 132.450 129.510 135.490 ;
        RECT 130.630 132.450 130.800 135.490 ;
        RECT 131.920 132.450 132.090 135.490 ;
        RECT 133.210 132.450 133.380 135.490 ;
        RECT 134.500 132.450 137.675 135.490 ;
        RECT 138.795 132.450 138.965 135.490 ;
        RECT 140.085 132.450 140.255 135.490 ;
        RECT 141.375 132.450 141.545 135.490 ;
        RECT 142.665 132.450 142.835 135.490 ;
        RECT 143.955 132.450 144.125 135.490 ;
        RECT 145.245 132.450 145.415 135.490 ;
        RECT 146.535 132.450 146.705 135.490 ;
        RECT 147.825 132.450 151.000 135.490 ;
        RECT 152.120 132.450 152.290 135.490 ;
        RECT 153.410 132.450 153.580 135.490 ;
        RECT 154.700 132.450 154.870 135.490 ;
        RECT 155.990 132.450 156.160 135.490 ;
        RECT 157.280 132.450 157.450 135.490 ;
        RECT 158.570 132.450 158.740 135.490 ;
        RECT 159.860 132.450 160.030 135.490 ;
        RECT 161.150 132.450 164.325 135.490 ;
        RECT 165.445 132.450 165.615 135.490 ;
        RECT 166.735 132.450 166.905 135.490 ;
        RECT 168.025 132.450 168.195 135.490 ;
        RECT 169.315 132.450 169.485 135.490 ;
        RECT 170.605 132.450 170.775 135.490 ;
        RECT 171.895 132.450 172.065 135.490 ;
        RECT 173.185 132.450 173.355 135.490 ;
        RECT 174.475 132.450 177.650 135.490 ;
        RECT 178.770 132.450 178.940 135.490 ;
        RECT 180.060 132.450 180.230 135.490 ;
        RECT 181.350 132.450 181.520 135.490 ;
        RECT 182.640 132.450 182.810 135.490 ;
        RECT 183.930 132.450 184.100 135.490 ;
        RECT 185.220 132.450 185.390 135.490 ;
        RECT 186.510 132.450 186.680 135.490 ;
        RECT 187.800 132.450 190.975 135.490 ;
        RECT 192.095 132.450 192.265 135.490 ;
        RECT 193.385 132.450 193.555 135.490 ;
        RECT 194.675 132.450 194.845 135.490 ;
        RECT 195.965 132.450 196.135 135.490 ;
        RECT 197.255 132.450 197.425 135.490 ;
        RECT 198.545 132.450 201.725 135.490 ;
        RECT 202.845 132.450 203.015 135.490 ;
        RECT 204.135 132.450 204.305 135.490 ;
        RECT 205.425 132.450 205.595 135.490 ;
        RECT 206.715 132.450 206.885 135.490 ;
        RECT 208.005 132.450 208.175 135.490 ;
        RECT 209.295 132.450 209.465 135.490 ;
        RECT 210.585 132.450 210.755 135.490 ;
        RECT 211.875 132.450 215.050 135.490 ;
        RECT 216.170 132.450 216.340 135.490 ;
        RECT 217.460 132.450 217.630 135.490 ;
        RECT 218.750 132.450 218.920 135.490 ;
        RECT 220.040 132.450 220.210 135.490 ;
        RECT 221.330 132.450 221.500 135.490 ;
        RECT 222.620 132.450 222.790 135.490 ;
        RECT 223.910 132.450 224.080 135.490 ;
        RECT 225.200 132.700 228.050 135.490 ;
        RECT 231.045 137.795 271.250 138.145 ;
        RECT 231.045 137.790 249.805 137.795 ;
        RECT 231.045 137.050 231.400 137.790 ;
        RECT 231.670 137.270 232.195 137.595 ;
        RECT 233.495 137.270 234.020 137.595 ;
        RECT 231.800 137.050 231.970 137.065 ;
        RECT 232.280 137.050 232.450 137.065 ;
        RECT 231.045 134.025 232.475 137.050 ;
        RECT 232.760 134.025 232.930 137.065 ;
        RECT 233.240 137.050 233.410 137.065 ;
        RECT 233.720 137.050 233.890 137.065 ;
        RECT 234.290 137.050 236.000 137.790 ;
        RECT 236.270 137.270 236.795 137.595 ;
        RECT 238.095 137.270 238.620 137.595 ;
        RECT 236.400 137.050 236.570 137.065 ;
        RECT 236.880 137.050 237.050 137.065 ;
        RECT 233.225 134.025 237.075 137.050 ;
        RECT 237.360 134.025 237.530 137.065 ;
        RECT 237.840 137.050 238.010 137.065 ;
        RECT 238.320 137.050 238.490 137.065 ;
        RECT 238.890 137.050 240.600 137.790 ;
        RECT 242.570 137.270 242.945 137.595 ;
        RECT 241.000 137.050 241.170 137.065 ;
        RECT 241.480 137.050 241.650 137.065 ;
        RECT 237.825 134.025 241.675 137.050 ;
        RECT 241.960 134.025 242.130 137.065 ;
        RECT 242.440 137.050 242.610 137.065 ;
        RECT 242.920 137.050 243.090 137.065 ;
        RECT 243.490 137.050 245.200 137.790 ;
        RECT 245.470 137.270 245.995 137.595 ;
        RECT 247.295 137.270 247.820 137.595 ;
        RECT 248.090 137.075 249.805 137.790 ;
        RECT 250.080 137.275 250.580 137.600 ;
        RECT 253.830 137.275 254.330 137.600 ;
        RECT 254.605 137.075 271.250 137.795 ;
        RECT 245.600 137.050 245.770 137.065 ;
        RECT 246.080 137.050 246.250 137.065 ;
        RECT 242.425 134.025 246.275 137.050 ;
        RECT 246.560 134.025 246.730 137.065 ;
        RECT 247.040 137.050 247.210 137.065 ;
        RECT 247.520 137.050 247.690 137.065 ;
        RECT 248.090 137.050 250.875 137.075 ;
        RECT 247.025 134.025 250.875 137.050 ;
        RECT 251.160 134.030 251.330 137.070 ;
        RECT 251.640 134.030 251.810 137.070 ;
        RECT 252.120 134.030 252.290 137.070 ;
        RECT 252.600 134.030 252.770 137.070 ;
        RECT 253.080 134.030 253.250 137.070 ;
        RECT 253.525 134.025 271.250 137.075 ;
        RECT 231.045 133.300 231.400 134.025 ;
        RECT 232.445 133.470 233.245 133.845 ;
        RECT 234.290 133.300 236.000 134.025 ;
        RECT 237.045 133.470 237.845 133.845 ;
        RECT 238.890 133.300 240.600 134.025 ;
        RECT 242.095 133.470 242.470 133.845 ;
        RECT 243.490 133.300 245.200 134.025 ;
        RECT 246.245 133.470 247.045 133.845 ;
        RECT 248.090 133.305 249.805 134.025 ;
        RECT 250.830 133.475 253.580 133.850 ;
        RECT 254.605 133.305 271.250 134.025 ;
        RECT 248.090 133.300 271.250 133.305 ;
        RECT 231.045 132.950 271.250 133.300 ;
        RECT 231.045 132.945 234.645 132.950 ;
        RECT 235.645 132.945 239.245 132.950 ;
        RECT 240.245 132.945 243.845 132.950 ;
        RECT 244.845 132.945 248.445 132.950 ;
        RECT 225.200 132.450 254.955 132.700 ;
        RECT 75.280 131.770 76.030 132.450 ;
        RECT 76.260 132.110 77.260 132.280 ;
        RECT 82.710 132.110 83.710 132.280 ;
        RECT 83.930 131.770 86.805 132.450 ;
        RECT 87.010 132.110 88.010 132.280 ;
        RECT 96.040 132.110 97.040 132.280 ;
        RECT 97.255 131.770 100.130 132.450 ;
        RECT 100.335 132.110 101.335 132.280 ;
        RECT 109.365 132.110 110.365 132.280 ;
        RECT 110.580 131.770 113.430 132.450 ;
        RECT 113.660 132.110 114.660 132.280 ;
        RECT 120.110 132.110 121.110 132.280 ;
        RECT 121.330 131.770 124.205 132.450 ;
        RECT 124.410 132.110 125.410 132.280 ;
        RECT 133.440 132.110 134.440 132.280 ;
        RECT 134.655 131.770 137.530 132.450 ;
        RECT 137.735 132.110 138.735 132.280 ;
        RECT 146.765 132.110 147.765 132.280 ;
        RECT 147.980 131.770 150.855 132.450 ;
        RECT 151.060 132.110 152.060 132.280 ;
        RECT 160.090 132.110 161.090 132.280 ;
        RECT 161.305 131.770 164.180 132.450 ;
        RECT 164.385 132.110 165.385 132.280 ;
        RECT 173.415 132.110 174.415 132.280 ;
        RECT 174.630 131.770 177.505 132.450 ;
        RECT 177.710 132.110 178.710 132.280 ;
        RECT 186.740 132.110 187.740 132.280 ;
        RECT 187.955 131.770 190.805 132.450 ;
        RECT 191.035 132.110 192.035 132.280 ;
        RECT 197.485 132.110 198.485 132.280 ;
        RECT 198.705 131.770 201.580 132.450 ;
        RECT 201.785 132.110 202.785 132.280 ;
        RECT 210.815 132.110 211.815 132.280 ;
        RECT 212.030 131.770 214.905 132.450 ;
        RECT 225.355 132.350 254.955 132.450 ;
        RECT 215.110 132.110 216.110 132.280 ;
        RECT 224.140 132.110 225.140 132.280 ;
        RECT 225.355 131.770 231.405 132.350 ;
        RECT 232.450 131.850 233.250 132.175 ;
        RECT 75.280 131.675 231.405 131.770 ;
        RECT 234.295 131.675 236.005 132.350 ;
        RECT 237.050 131.850 237.850 132.175 ;
        RECT 238.895 131.675 240.605 132.350 ;
        RECT 242.100 131.850 242.475 132.175 ;
        RECT 243.495 131.675 245.205 132.350 ;
        RECT 246.250 131.850 247.050 132.175 ;
        RECT 248.095 131.675 249.805 132.350 ;
        RECT 250.830 131.850 253.580 132.175 ;
        RECT 254.605 131.675 254.955 132.350 ;
        RECT 75.280 130.625 232.475 131.675 ;
        RECT 232.765 130.630 232.935 131.670 ;
        RECT 233.225 130.625 237.075 131.675 ;
        RECT 237.365 130.630 237.535 131.670 ;
        RECT 237.825 130.625 241.675 131.675 ;
        RECT 241.965 130.630 242.135 131.670 ;
        RECT 242.425 130.625 246.275 131.675 ;
        RECT 246.565 130.630 246.735 131.670 ;
        RECT 247.025 130.625 250.875 131.675 ;
        RECT 251.160 130.630 251.330 131.670 ;
        RECT 251.640 130.630 251.810 131.670 ;
        RECT 252.120 130.630 252.290 131.670 ;
        RECT 252.600 130.630 252.770 131.670 ;
        RECT 253.080 130.630 253.250 131.670 ;
        RECT 253.525 130.625 254.955 131.675 ;
        RECT 75.280 129.950 231.405 130.625 ;
        RECT 231.675 130.125 232.200 130.450 ;
        RECT 233.500 130.125 234.025 130.450 ;
        RECT 234.295 129.950 236.005 130.625 ;
        RECT 236.275 130.125 236.800 130.450 ;
        RECT 238.100 130.125 238.625 130.450 ;
        RECT 238.895 129.950 240.605 130.625 ;
        RECT 242.575 130.125 242.950 130.450 ;
        RECT 243.495 129.950 245.205 130.625 ;
        RECT 245.475 130.125 246.000 130.450 ;
        RECT 247.300 130.125 247.825 130.450 ;
        RECT 248.095 129.950 249.805 130.625 ;
        RECT 250.080 130.125 250.580 130.450 ;
        RECT 253.830 130.125 254.330 130.450 ;
        RECT 254.605 129.950 254.955 130.625 ;
        RECT 75.280 129.600 254.955 129.950 ;
        RECT 256.625 132.090 271.250 132.950 ;
        RECT 75.280 129.445 228.050 129.600 ;
        RECT 97.130 128.800 212.490 128.815 ;
        RECT 75.275 128.645 212.675 128.800 ;
        RECT 75.275 121.525 97.300 128.645 ;
        RECT 97.780 126.005 98.130 128.165 ;
        RECT 98.610 126.005 98.960 128.165 ;
        RECT 99.440 126.005 99.790 128.165 ;
        RECT 100.270 126.005 100.620 128.165 ;
        RECT 101.100 126.005 101.450 128.165 ;
        RECT 101.930 126.005 102.280 128.165 ;
        RECT 102.760 126.005 103.110 128.165 ;
        RECT 103.590 126.005 103.940 128.165 ;
        RECT 104.420 126.005 104.770 128.165 ;
        RECT 105.250 126.005 105.600 128.165 ;
        RECT 106.080 126.005 106.430 128.165 ;
        RECT 106.910 126.005 107.260 128.165 ;
        RECT 107.740 126.005 108.090 128.165 ;
        RECT 108.570 126.005 108.920 128.165 ;
        RECT 109.400 126.005 109.750 128.165 ;
        RECT 110.230 126.005 110.580 128.165 ;
        RECT 111.060 126.005 111.410 128.165 ;
        RECT 111.890 126.005 112.240 128.165 ;
        RECT 112.720 126.005 113.070 128.165 ;
        RECT 113.550 126.005 113.900 128.165 ;
        RECT 114.380 126.005 114.730 128.165 ;
        RECT 115.210 126.005 115.560 128.165 ;
        RECT 116.040 126.005 116.390 128.165 ;
        RECT 116.870 126.005 117.220 128.165 ;
        RECT 117.700 126.005 118.050 128.165 ;
        RECT 118.530 126.005 118.880 128.165 ;
        RECT 119.360 126.005 119.710 128.165 ;
        RECT 120.190 126.005 120.540 128.165 ;
        RECT 121.020 126.005 121.370 128.165 ;
        RECT 121.850 126.005 122.200 128.165 ;
        RECT 122.680 126.005 123.030 128.165 ;
        RECT 123.510 126.005 123.860 128.165 ;
        RECT 124.340 126.005 124.690 128.165 ;
        RECT 125.170 126.005 125.520 128.165 ;
        RECT 126.000 126.005 126.350 128.165 ;
        RECT 126.830 126.005 127.180 128.165 ;
        RECT 127.660 126.005 128.010 128.165 ;
        RECT 128.490 126.005 128.840 128.165 ;
        RECT 129.320 126.005 129.670 128.165 ;
        RECT 130.150 126.005 130.500 128.165 ;
        RECT 130.980 126.005 131.330 128.165 ;
        RECT 131.810 126.005 132.160 128.165 ;
        RECT 132.640 126.005 132.990 128.165 ;
        RECT 133.470 126.005 133.820 128.165 ;
        RECT 134.300 126.005 134.650 128.165 ;
        RECT 135.130 126.005 135.480 128.165 ;
        RECT 135.960 126.005 136.310 128.165 ;
        RECT 136.790 126.005 137.140 128.165 ;
        RECT 137.620 126.005 137.970 128.165 ;
        RECT 138.450 126.005 138.800 128.165 ;
        RECT 139.280 126.005 139.630 128.165 ;
        RECT 140.110 126.005 140.460 128.165 ;
        RECT 140.940 126.005 141.290 128.165 ;
        RECT 141.770 126.005 142.120 128.165 ;
        RECT 142.600 126.005 142.950 128.165 ;
        RECT 143.430 126.005 143.780 128.165 ;
        RECT 144.260 126.005 144.610 128.165 ;
        RECT 145.090 126.005 145.440 128.165 ;
        RECT 145.920 126.005 146.270 128.165 ;
        RECT 146.750 126.005 147.100 128.165 ;
        RECT 147.580 126.005 147.930 128.165 ;
        RECT 148.410 126.005 148.760 128.165 ;
        RECT 149.240 126.005 149.590 128.165 ;
        RECT 150.070 126.005 150.420 128.165 ;
        RECT 150.900 126.005 151.250 128.165 ;
        RECT 151.730 126.005 152.080 128.165 ;
        RECT 152.560 126.005 152.910 128.165 ;
        RECT 153.390 126.005 153.740 128.165 ;
        RECT 154.220 126.005 154.570 128.165 ;
        RECT 155.050 126.005 155.400 128.165 ;
        RECT 155.880 126.005 156.230 128.165 ;
        RECT 156.710 126.005 157.060 128.165 ;
        RECT 157.540 126.005 157.890 128.165 ;
        RECT 158.370 126.005 158.720 128.165 ;
        RECT 159.200 126.005 159.550 128.165 ;
        RECT 160.030 126.005 160.380 128.165 ;
        RECT 160.860 126.005 161.210 128.165 ;
        RECT 161.690 126.005 162.040 128.165 ;
        RECT 162.520 126.005 162.870 128.165 ;
        RECT 163.350 126.005 163.700 128.165 ;
        RECT 164.180 126.005 164.530 128.165 ;
        RECT 165.010 126.005 165.360 128.165 ;
        RECT 165.840 126.005 166.190 128.165 ;
        RECT 166.670 126.005 167.020 128.165 ;
        RECT 167.500 126.005 167.850 128.165 ;
        RECT 168.330 126.005 168.680 128.165 ;
        RECT 169.160 126.005 169.510 128.165 ;
        RECT 169.990 126.005 170.340 128.165 ;
        RECT 170.820 126.005 171.170 128.165 ;
        RECT 171.650 126.005 172.000 128.165 ;
        RECT 172.480 126.005 172.830 128.165 ;
        RECT 173.310 126.005 173.660 128.165 ;
        RECT 174.140 126.005 174.490 128.165 ;
        RECT 174.970 126.005 175.320 128.165 ;
        RECT 175.800 126.005 176.150 128.165 ;
        RECT 176.630 126.005 176.980 128.165 ;
        RECT 177.460 126.005 177.810 128.165 ;
        RECT 178.290 126.005 178.640 128.165 ;
        RECT 179.120 126.005 179.470 128.165 ;
        RECT 179.950 126.005 180.300 128.165 ;
        RECT 180.780 126.005 181.130 128.165 ;
        RECT 181.610 126.005 181.960 128.165 ;
        RECT 182.440 126.005 182.790 128.165 ;
        RECT 183.270 126.005 183.620 128.165 ;
        RECT 184.100 126.005 184.450 128.165 ;
        RECT 184.930 126.005 185.280 128.165 ;
        RECT 185.760 126.005 186.110 128.165 ;
        RECT 186.590 126.005 186.940 128.165 ;
        RECT 187.420 126.005 187.770 128.165 ;
        RECT 188.250 126.005 188.600 128.165 ;
        RECT 189.080 126.005 189.430 128.165 ;
        RECT 189.910 126.005 190.260 128.165 ;
        RECT 190.740 126.005 191.090 128.165 ;
        RECT 191.570 126.005 191.920 128.165 ;
        RECT 192.400 126.005 192.750 128.165 ;
        RECT 193.230 126.005 193.580 128.165 ;
        RECT 194.060 126.005 194.410 128.165 ;
        RECT 194.890 126.005 195.240 128.165 ;
        RECT 195.720 126.005 196.070 128.165 ;
        RECT 196.550 126.005 196.900 128.165 ;
        RECT 197.380 126.005 197.730 128.165 ;
        RECT 198.210 126.005 198.560 128.165 ;
        RECT 199.040 126.005 199.390 128.165 ;
        RECT 199.870 126.005 200.220 128.165 ;
        RECT 200.700 126.005 201.050 128.165 ;
        RECT 201.530 126.005 201.880 128.165 ;
        RECT 202.360 126.005 202.710 128.165 ;
        RECT 203.190 126.005 203.540 128.165 ;
        RECT 204.020 126.005 204.370 128.165 ;
        RECT 204.850 126.005 205.200 128.165 ;
        RECT 205.680 126.005 206.030 128.165 ;
        RECT 206.510 126.005 206.860 128.165 ;
        RECT 207.340 126.005 207.690 128.165 ;
        RECT 208.170 126.005 208.520 128.165 ;
        RECT 209.000 126.005 209.350 128.165 ;
        RECT 209.830 126.005 210.180 128.165 ;
        RECT 210.660 126.005 211.010 128.165 ;
        RECT 211.490 126.005 211.840 128.165 ;
        RECT 212.320 125.400 212.675 128.645 ;
        RECT 215.625 125.400 228.050 129.445 ;
        RECT 97.780 122.005 98.130 124.165 ;
        RECT 98.610 122.005 98.960 124.165 ;
        RECT 99.440 122.005 99.790 124.165 ;
        RECT 100.270 122.005 100.620 124.165 ;
        RECT 101.100 122.005 101.450 124.165 ;
        RECT 101.930 122.005 102.280 124.165 ;
        RECT 102.760 122.005 103.110 124.165 ;
        RECT 103.590 122.005 103.940 124.165 ;
        RECT 104.420 122.005 104.770 124.165 ;
        RECT 105.250 122.005 105.600 124.165 ;
        RECT 106.080 122.005 106.430 124.165 ;
        RECT 106.910 122.005 107.260 124.165 ;
        RECT 107.740 122.005 108.090 124.165 ;
        RECT 108.570 122.005 108.920 124.165 ;
        RECT 109.400 122.005 109.750 124.165 ;
        RECT 110.230 122.005 110.580 124.165 ;
        RECT 111.060 122.005 111.410 124.165 ;
        RECT 111.890 122.005 112.240 124.165 ;
        RECT 112.720 122.005 113.070 124.165 ;
        RECT 113.550 122.005 113.900 124.165 ;
        RECT 114.380 122.005 114.730 124.165 ;
        RECT 115.210 122.005 115.560 124.165 ;
        RECT 116.040 122.005 116.390 124.165 ;
        RECT 116.870 122.005 117.220 124.165 ;
        RECT 117.700 122.005 118.050 124.165 ;
        RECT 118.530 122.005 118.880 124.165 ;
        RECT 119.360 122.005 119.710 124.165 ;
        RECT 120.190 122.005 120.540 124.165 ;
        RECT 121.020 122.005 121.370 124.165 ;
        RECT 121.850 122.005 122.200 124.165 ;
        RECT 122.680 122.005 123.030 124.165 ;
        RECT 123.510 122.005 123.860 124.165 ;
        RECT 124.340 122.005 124.690 124.165 ;
        RECT 125.170 122.005 125.520 124.165 ;
        RECT 126.000 122.005 126.350 124.165 ;
        RECT 126.830 122.005 127.180 124.165 ;
        RECT 127.660 122.005 128.010 124.165 ;
        RECT 128.490 122.005 128.840 124.165 ;
        RECT 129.320 122.005 129.670 124.165 ;
        RECT 130.150 122.005 130.500 124.165 ;
        RECT 130.980 122.005 131.330 124.165 ;
        RECT 131.810 122.005 132.160 124.165 ;
        RECT 132.640 122.005 132.990 124.165 ;
        RECT 133.470 122.005 133.820 124.165 ;
        RECT 134.300 122.005 134.650 124.165 ;
        RECT 135.130 122.005 135.480 124.165 ;
        RECT 135.960 122.005 136.310 124.165 ;
        RECT 136.790 122.005 137.140 124.165 ;
        RECT 137.620 122.005 137.970 124.165 ;
        RECT 138.450 122.005 138.800 124.165 ;
        RECT 139.280 122.005 139.630 124.165 ;
        RECT 140.110 122.005 140.460 124.165 ;
        RECT 140.940 122.005 141.290 124.165 ;
        RECT 141.770 122.005 142.120 124.165 ;
        RECT 142.600 122.005 142.950 124.165 ;
        RECT 143.430 122.005 143.780 124.165 ;
        RECT 144.260 122.005 144.610 124.165 ;
        RECT 145.090 122.005 145.440 124.165 ;
        RECT 145.920 122.005 146.270 124.165 ;
        RECT 146.750 122.005 147.100 124.165 ;
        RECT 147.580 122.005 147.930 124.165 ;
        RECT 148.410 122.005 148.760 124.165 ;
        RECT 149.240 122.005 149.590 124.165 ;
        RECT 150.070 122.005 150.420 124.165 ;
        RECT 150.900 122.005 151.250 124.165 ;
        RECT 151.730 122.005 152.080 124.165 ;
        RECT 152.560 122.005 152.910 124.165 ;
        RECT 153.390 122.005 153.740 124.165 ;
        RECT 154.220 122.005 154.570 124.165 ;
        RECT 155.050 122.005 155.400 124.165 ;
        RECT 155.880 122.005 156.230 124.165 ;
        RECT 156.710 122.005 157.060 124.165 ;
        RECT 157.540 122.005 157.890 124.165 ;
        RECT 158.370 122.005 158.720 124.165 ;
        RECT 159.200 122.005 159.550 124.165 ;
        RECT 160.030 122.005 160.380 124.165 ;
        RECT 160.860 122.005 161.210 124.165 ;
        RECT 161.690 122.005 162.040 124.165 ;
        RECT 162.520 122.005 162.870 124.165 ;
        RECT 163.350 122.005 163.700 124.165 ;
        RECT 164.180 122.005 164.530 124.165 ;
        RECT 165.010 122.005 165.360 124.165 ;
        RECT 165.840 122.005 166.190 124.165 ;
        RECT 166.670 122.005 167.020 124.165 ;
        RECT 167.500 122.005 167.850 124.165 ;
        RECT 168.330 122.005 168.680 124.165 ;
        RECT 169.160 122.005 169.510 124.165 ;
        RECT 169.990 122.005 170.340 124.165 ;
        RECT 170.820 122.005 171.170 124.165 ;
        RECT 171.650 122.005 172.000 124.165 ;
        RECT 172.480 122.005 172.830 124.165 ;
        RECT 173.310 122.005 173.660 124.165 ;
        RECT 174.140 122.005 174.490 124.165 ;
        RECT 174.970 122.005 175.320 124.165 ;
        RECT 175.800 122.005 176.150 124.165 ;
        RECT 176.630 122.005 176.980 124.165 ;
        RECT 177.460 122.005 177.810 124.165 ;
        RECT 178.290 122.005 178.640 124.165 ;
        RECT 179.120 122.005 179.470 124.165 ;
        RECT 179.950 122.005 180.300 124.165 ;
        RECT 180.780 122.005 181.130 124.165 ;
        RECT 181.610 122.005 181.960 124.165 ;
        RECT 182.440 122.005 182.790 124.165 ;
        RECT 183.270 122.005 183.620 124.165 ;
        RECT 184.100 122.005 184.450 124.165 ;
        RECT 184.930 122.005 185.280 124.165 ;
        RECT 185.760 122.005 186.110 124.165 ;
        RECT 186.590 122.005 186.940 124.165 ;
        RECT 187.420 122.005 187.770 124.165 ;
        RECT 188.250 122.005 188.600 124.165 ;
        RECT 189.080 122.005 189.430 124.165 ;
        RECT 189.910 122.005 190.260 124.165 ;
        RECT 190.740 122.005 191.090 124.165 ;
        RECT 191.570 122.005 191.920 124.165 ;
        RECT 192.400 122.005 192.750 124.165 ;
        RECT 193.230 122.005 193.580 124.165 ;
        RECT 194.060 122.005 194.410 124.165 ;
        RECT 194.890 122.005 195.240 124.165 ;
        RECT 195.720 122.005 196.070 124.165 ;
        RECT 196.550 122.005 196.900 124.165 ;
        RECT 197.380 122.005 197.730 124.165 ;
        RECT 198.210 122.005 198.560 124.165 ;
        RECT 199.040 122.005 199.390 124.165 ;
        RECT 199.870 122.005 200.220 124.165 ;
        RECT 200.700 122.005 201.050 124.165 ;
        RECT 201.530 122.005 201.880 124.165 ;
        RECT 202.360 122.005 202.710 124.165 ;
        RECT 203.190 122.005 203.540 124.165 ;
        RECT 204.020 122.005 204.370 124.165 ;
        RECT 204.850 122.005 205.200 124.165 ;
        RECT 205.680 122.005 206.030 124.165 ;
        RECT 206.510 122.005 206.860 124.165 ;
        RECT 207.340 122.005 207.690 124.165 ;
        RECT 208.170 122.005 208.520 124.165 ;
        RECT 209.000 122.005 209.350 124.165 ;
        RECT 209.830 122.005 210.180 124.165 ;
        RECT 210.660 122.005 211.010 124.165 ;
        RECT 211.490 122.005 211.840 124.165 ;
        RECT 212.320 123.400 228.050 125.400 ;
        RECT 231.050 128.850 233.700 128.855 ;
        RECT 231.050 128.500 254.955 128.850 ;
        RECT 231.050 124.010 231.425 128.500 ;
        RECT 233.325 128.495 254.955 128.500 ;
        RECT 233.325 128.490 249.805 128.495 ;
        RECT 231.950 127.955 232.800 128.330 ;
        RECT 231.810 124.735 231.980 127.775 ;
        RECT 232.290 124.735 232.460 127.775 ;
        RECT 232.770 124.735 232.940 127.775 ;
        RECT 233.325 127.750 236.000 128.490 ;
        RECT 236.270 127.970 236.795 128.295 ;
        RECT 238.095 127.970 238.620 128.295 ;
        RECT 236.400 127.750 236.570 127.765 ;
        RECT 236.880 127.750 237.050 127.765 ;
        RECT 233.325 124.725 237.075 127.750 ;
        RECT 237.360 124.725 237.530 127.765 ;
        RECT 237.840 127.750 238.010 127.765 ;
        RECT 238.320 127.750 238.490 127.765 ;
        RECT 238.890 127.750 240.600 128.490 ;
        RECT 242.570 127.970 242.945 128.295 ;
        RECT 241.000 127.750 241.170 127.765 ;
        RECT 241.480 127.750 241.650 127.765 ;
        RECT 237.825 124.725 241.675 127.750 ;
        RECT 241.960 124.725 242.130 127.765 ;
        RECT 242.440 127.750 242.610 127.765 ;
        RECT 242.920 127.750 243.090 127.765 ;
        RECT 243.490 127.750 245.200 128.490 ;
        RECT 245.470 127.970 245.995 128.295 ;
        RECT 247.295 127.970 247.820 128.295 ;
        RECT 248.090 127.775 249.805 128.490 ;
        RECT 250.080 127.975 250.580 128.300 ;
        RECT 253.830 127.975 254.330 128.300 ;
        RECT 254.605 127.775 254.955 128.495 ;
        RECT 245.600 127.750 245.770 127.765 ;
        RECT 246.080 127.750 246.250 127.765 ;
        RECT 242.425 124.725 246.275 127.750 ;
        RECT 246.560 124.725 246.730 127.765 ;
        RECT 247.040 127.750 247.210 127.765 ;
        RECT 247.520 127.750 247.690 127.765 ;
        RECT 248.090 127.750 250.875 127.775 ;
        RECT 247.025 124.725 250.875 127.750 ;
        RECT 251.160 124.730 251.330 127.770 ;
        RECT 251.640 124.730 251.810 127.770 ;
        RECT 252.120 124.730 252.290 127.770 ;
        RECT 252.600 124.730 252.770 127.770 ;
        RECT 253.080 124.730 253.250 127.770 ;
        RECT 253.525 124.725 254.955 127.775 ;
        RECT 256.625 127.600 256.975 132.090 ;
        RECT 257.540 131.545 259.290 131.920 ;
        RECT 268.590 131.545 270.340 131.920 ;
        RECT 257.375 128.325 257.545 131.365 ;
        RECT 257.855 128.325 258.025 131.365 ;
        RECT 258.335 128.325 258.505 131.365 ;
        RECT 258.815 128.325 258.985 131.365 ;
        RECT 259.295 128.325 259.465 131.365 ;
        RECT 259.775 128.325 259.945 131.365 ;
        RECT 260.255 128.325 260.425 131.365 ;
        RECT 260.735 128.325 260.905 131.365 ;
        RECT 261.215 128.325 261.385 131.365 ;
        RECT 261.695 128.325 261.865 131.365 ;
        RECT 262.175 128.325 262.345 131.365 ;
        RECT 262.655 128.325 262.825 131.365 ;
        RECT 263.135 128.325 263.305 131.365 ;
        RECT 263.615 128.325 263.785 131.365 ;
        RECT 264.095 128.325 264.265 131.365 ;
        RECT 264.575 128.325 264.745 131.365 ;
        RECT 265.055 128.325 265.225 131.365 ;
        RECT 265.535 128.325 265.705 131.365 ;
        RECT 266.015 128.325 266.185 131.365 ;
        RECT 266.495 128.325 266.665 131.365 ;
        RECT 266.975 128.325 267.145 131.365 ;
        RECT 267.455 128.325 267.625 131.365 ;
        RECT 267.935 128.325 268.105 131.365 ;
        RECT 268.415 128.325 268.585 131.365 ;
        RECT 268.895 128.325 269.065 131.365 ;
        RECT 269.375 128.325 269.545 131.365 ;
        RECT 269.855 128.325 270.025 131.365 ;
        RECT 270.335 128.325 270.505 131.365 ;
        RECT 259.465 127.770 268.415 128.145 ;
        RECT 270.900 127.600 271.250 132.090 ;
        RECT 256.625 127.250 271.250 127.600 ;
        RECT 233.325 124.010 236.000 124.725 ;
        RECT 237.045 124.170 237.845 124.545 ;
        RECT 231.050 124.000 236.000 124.010 ;
        RECT 238.890 124.000 240.600 124.725 ;
        RECT 242.095 124.170 242.470 124.545 ;
        RECT 243.490 124.000 245.200 124.725 ;
        RECT 246.245 124.170 247.045 124.545 ;
        RECT 248.090 124.005 249.805 124.725 ;
        RECT 250.830 124.175 253.580 124.550 ;
        RECT 254.605 124.005 254.955 124.725 ;
        RECT 248.090 124.000 254.955 124.005 ;
        RECT 231.050 123.655 254.955 124.000 ;
        RECT 233.325 123.650 254.955 123.655 ;
        RECT 256.625 126.650 271.250 127.000 ;
        RECT 256.625 124.250 256.975 126.650 ;
        RECT 257.540 126.150 259.290 126.475 ;
        RECT 268.590 126.150 270.340 126.475 ;
        RECT 257.375 124.930 257.545 125.970 ;
        RECT 257.855 124.930 258.025 125.970 ;
        RECT 258.335 124.930 258.505 125.970 ;
        RECT 258.815 124.930 258.985 125.970 ;
        RECT 259.295 124.930 259.465 125.970 ;
        RECT 259.775 124.930 259.945 125.970 ;
        RECT 260.255 124.930 260.425 125.970 ;
        RECT 260.735 124.930 260.905 125.970 ;
        RECT 261.215 124.930 261.385 125.970 ;
        RECT 261.695 124.930 261.865 125.970 ;
        RECT 262.175 124.930 262.345 125.970 ;
        RECT 262.655 124.930 262.825 125.970 ;
        RECT 263.135 124.930 263.305 125.970 ;
        RECT 263.615 124.930 263.785 125.970 ;
        RECT 264.095 124.930 264.265 125.970 ;
        RECT 264.575 124.930 264.745 125.970 ;
        RECT 265.055 124.930 265.225 125.970 ;
        RECT 265.535 124.930 265.705 125.970 ;
        RECT 266.015 124.930 266.185 125.970 ;
        RECT 266.495 124.930 266.665 125.970 ;
        RECT 266.975 124.930 267.145 125.970 ;
        RECT 267.455 124.930 267.625 125.970 ;
        RECT 267.935 124.930 268.105 125.970 ;
        RECT 268.415 124.930 268.585 125.970 ;
        RECT 268.895 124.930 269.065 125.970 ;
        RECT 269.375 124.930 269.545 125.970 ;
        RECT 269.855 124.930 270.025 125.970 ;
        RECT 270.335 124.930 270.505 125.970 ;
        RECT 259.465 124.425 268.415 124.750 ;
        RECT 270.900 124.250 271.250 126.650 ;
        RECT 235.645 123.645 239.245 123.650 ;
        RECT 240.245 123.645 243.845 123.650 ;
        RECT 244.845 123.645 248.445 123.650 ;
        RECT 212.320 123.375 254.955 123.400 ;
        RECT 256.625 123.375 271.250 124.250 ;
        RECT 212.320 123.050 271.250 123.375 ;
        RECT 212.320 121.525 231.425 123.050 ;
        RECT 233.325 122.375 236.005 123.050 ;
        RECT 237.050 122.550 237.850 122.875 ;
        RECT 238.895 122.375 240.605 123.050 ;
        RECT 242.100 122.550 242.475 122.875 ;
        RECT 243.495 122.375 245.205 123.050 ;
        RECT 246.250 122.550 247.050 122.875 ;
        RECT 248.095 122.375 249.805 123.050 ;
        RECT 250.830 122.550 253.580 122.875 ;
        RECT 254.605 122.375 271.250 123.050 ;
        RECT 75.275 120.650 231.425 121.525 ;
        RECT 231.810 121.330 231.980 122.370 ;
        RECT 232.290 121.330 232.460 122.370 ;
        RECT 232.770 121.330 232.940 122.370 ;
        RECT 233.325 121.325 237.075 122.375 ;
        RECT 237.365 121.330 237.535 122.370 ;
        RECT 237.825 121.325 241.675 122.375 ;
        RECT 241.965 121.330 242.135 122.370 ;
        RECT 242.425 121.325 246.275 122.375 ;
        RECT 246.565 121.330 246.735 122.370 ;
        RECT 247.025 121.325 250.875 122.375 ;
        RECT 251.160 121.330 251.330 122.370 ;
        RECT 251.640 121.330 251.810 122.370 ;
        RECT 252.120 121.330 252.290 122.370 ;
        RECT 252.600 121.330 252.770 122.370 ;
        RECT 253.080 121.330 253.250 122.370 ;
        RECT 253.525 121.325 271.250 122.375 ;
        RECT 231.950 120.825 232.800 121.150 ;
        RECT 233.325 120.650 236.005 121.325 ;
        RECT 236.275 120.825 236.800 121.150 ;
        RECT 238.100 120.825 238.625 121.150 ;
        RECT 238.895 120.650 240.605 121.325 ;
        RECT 242.575 120.825 242.950 121.150 ;
        RECT 243.495 120.650 245.205 121.325 ;
        RECT 245.475 120.825 246.000 121.150 ;
        RECT 247.300 120.825 247.825 121.150 ;
        RECT 248.095 120.650 249.805 121.325 ;
        RECT 250.080 120.825 250.580 121.150 ;
        RECT 253.830 120.825 254.330 121.150 ;
        RECT 254.605 120.650 271.250 121.325 ;
        RECT 75.275 119.450 271.250 120.650 ;
        RECT 75.275 104.370 228.050 119.450 ;
        RECT 231.050 115.025 271.250 119.450 ;
        RECT 231.050 105.495 271.250 110.775 ;
        RECT 75.275 97.250 97.300 104.370 ;
        RECT 97.780 101.730 98.130 103.890 ;
        RECT 98.610 101.730 98.960 103.890 ;
        RECT 99.440 101.730 99.790 103.890 ;
        RECT 100.270 101.730 100.620 103.890 ;
        RECT 101.100 101.730 101.450 103.890 ;
        RECT 101.930 101.730 102.280 103.890 ;
        RECT 102.760 101.730 103.110 103.890 ;
        RECT 103.590 101.730 103.940 103.890 ;
        RECT 104.420 101.730 104.770 103.890 ;
        RECT 105.250 101.730 105.600 103.890 ;
        RECT 106.080 101.730 106.430 103.890 ;
        RECT 106.910 101.730 107.260 103.890 ;
        RECT 107.740 101.730 108.090 103.890 ;
        RECT 108.570 101.730 108.920 103.890 ;
        RECT 109.400 101.730 109.750 103.890 ;
        RECT 110.230 101.730 110.580 103.890 ;
        RECT 111.060 101.730 111.410 103.890 ;
        RECT 111.890 101.730 112.240 103.890 ;
        RECT 112.720 101.730 113.070 103.890 ;
        RECT 113.550 101.730 113.900 103.890 ;
        RECT 114.380 101.730 114.730 103.890 ;
        RECT 115.210 101.730 115.560 103.890 ;
        RECT 116.040 101.730 116.390 103.890 ;
        RECT 116.870 101.730 117.220 103.890 ;
        RECT 117.700 101.730 118.050 103.890 ;
        RECT 118.530 101.730 118.880 103.890 ;
        RECT 119.360 101.730 119.710 103.890 ;
        RECT 120.190 101.730 120.540 103.890 ;
        RECT 121.020 101.730 121.370 103.890 ;
        RECT 121.850 101.730 122.200 103.890 ;
        RECT 122.680 101.730 123.030 103.890 ;
        RECT 123.510 101.730 123.860 103.890 ;
        RECT 124.340 101.730 124.690 103.890 ;
        RECT 125.170 101.730 125.520 103.890 ;
        RECT 126.000 101.730 126.350 103.890 ;
        RECT 126.830 101.730 127.180 103.890 ;
        RECT 127.660 101.730 128.010 103.890 ;
        RECT 128.490 101.730 128.840 103.890 ;
        RECT 129.320 101.730 129.670 103.890 ;
        RECT 130.150 101.730 130.500 103.890 ;
        RECT 130.980 101.730 131.330 103.890 ;
        RECT 131.810 101.730 132.160 103.890 ;
        RECT 132.640 101.730 132.990 103.890 ;
        RECT 133.470 101.730 133.820 103.890 ;
        RECT 134.300 101.730 134.650 103.890 ;
        RECT 135.130 101.730 135.480 103.890 ;
        RECT 135.960 101.730 136.310 103.890 ;
        RECT 136.790 101.730 137.140 103.890 ;
        RECT 137.620 101.730 137.970 103.890 ;
        RECT 138.450 101.730 138.800 103.890 ;
        RECT 139.280 101.730 139.630 103.890 ;
        RECT 140.110 101.730 140.460 103.890 ;
        RECT 140.940 101.730 141.290 103.890 ;
        RECT 141.770 101.730 142.120 103.890 ;
        RECT 142.600 101.730 142.950 103.890 ;
        RECT 143.430 101.730 143.780 103.890 ;
        RECT 144.260 101.730 144.610 103.890 ;
        RECT 145.090 101.730 145.440 103.890 ;
        RECT 145.920 101.730 146.270 103.890 ;
        RECT 146.750 101.730 147.100 103.890 ;
        RECT 147.580 101.730 147.930 103.890 ;
        RECT 148.410 101.730 148.760 103.890 ;
        RECT 149.240 101.730 149.590 103.890 ;
        RECT 150.070 101.730 150.420 103.890 ;
        RECT 150.900 101.730 151.250 103.890 ;
        RECT 151.730 101.730 152.080 103.890 ;
        RECT 152.560 101.730 152.910 103.890 ;
        RECT 153.390 101.730 153.740 103.890 ;
        RECT 154.220 101.730 154.570 103.890 ;
        RECT 155.050 101.730 155.400 103.890 ;
        RECT 155.880 101.730 156.230 103.890 ;
        RECT 156.710 101.730 157.060 103.890 ;
        RECT 157.540 101.730 157.890 103.890 ;
        RECT 158.370 101.730 158.720 103.890 ;
        RECT 159.200 101.730 159.550 103.890 ;
        RECT 160.030 101.730 160.380 103.890 ;
        RECT 160.860 101.730 161.210 103.890 ;
        RECT 161.690 101.730 162.040 103.890 ;
        RECT 162.520 101.730 162.870 103.890 ;
        RECT 163.350 101.730 163.700 103.890 ;
        RECT 164.180 101.730 164.530 103.890 ;
        RECT 165.010 101.730 165.360 103.890 ;
        RECT 165.840 101.730 166.190 103.890 ;
        RECT 166.670 101.730 167.020 103.890 ;
        RECT 167.500 101.730 167.850 103.890 ;
        RECT 168.330 101.730 168.680 103.890 ;
        RECT 169.160 101.730 169.510 103.890 ;
        RECT 169.990 101.730 170.340 103.890 ;
        RECT 170.820 101.730 171.170 103.890 ;
        RECT 171.650 101.730 172.000 103.890 ;
        RECT 172.480 101.730 172.830 103.890 ;
        RECT 173.310 101.730 173.660 103.890 ;
        RECT 174.140 101.730 174.490 103.890 ;
        RECT 174.970 101.730 175.320 103.890 ;
        RECT 175.800 101.730 176.150 103.890 ;
        RECT 176.630 101.730 176.980 103.890 ;
        RECT 177.460 101.730 177.810 103.890 ;
        RECT 178.290 101.730 178.640 103.890 ;
        RECT 179.120 101.730 179.470 103.890 ;
        RECT 179.950 101.730 180.300 103.890 ;
        RECT 180.780 101.730 181.130 103.890 ;
        RECT 181.610 101.730 181.960 103.890 ;
        RECT 182.440 101.730 182.790 103.890 ;
        RECT 183.270 101.730 183.620 103.890 ;
        RECT 184.100 101.730 184.450 103.890 ;
        RECT 184.930 101.730 185.280 103.890 ;
        RECT 185.760 101.730 186.110 103.890 ;
        RECT 186.590 101.730 186.940 103.890 ;
        RECT 187.420 101.730 187.770 103.890 ;
        RECT 188.250 101.730 188.600 103.890 ;
        RECT 189.080 101.730 189.430 103.890 ;
        RECT 189.910 101.730 190.260 103.890 ;
        RECT 190.740 101.730 191.090 103.890 ;
        RECT 191.570 101.730 191.920 103.890 ;
        RECT 192.400 101.730 192.750 103.890 ;
        RECT 193.230 101.730 193.580 103.890 ;
        RECT 194.060 101.730 194.410 103.890 ;
        RECT 194.890 101.730 195.240 103.890 ;
        RECT 195.720 101.730 196.070 103.890 ;
        RECT 196.550 101.730 196.900 103.890 ;
        RECT 197.380 101.730 197.730 103.890 ;
        RECT 198.210 101.730 198.560 103.890 ;
        RECT 199.040 101.730 199.390 103.890 ;
        RECT 199.870 101.730 200.220 103.890 ;
        RECT 200.700 101.730 201.050 103.890 ;
        RECT 201.530 101.730 201.880 103.890 ;
        RECT 202.360 101.730 202.710 103.890 ;
        RECT 203.190 101.730 203.540 103.890 ;
        RECT 204.020 101.730 204.370 103.890 ;
        RECT 204.850 101.730 205.200 103.890 ;
        RECT 205.680 101.730 206.030 103.890 ;
        RECT 206.510 101.730 206.860 103.890 ;
        RECT 207.340 101.730 207.690 103.890 ;
        RECT 208.170 101.730 208.520 103.890 ;
        RECT 209.000 101.730 209.350 103.890 ;
        RECT 209.830 101.730 210.180 103.890 ;
        RECT 210.660 101.730 211.010 103.890 ;
        RECT 211.490 101.730 211.840 103.890 ;
        RECT 212.320 100.500 228.050 104.370 ;
        RECT 97.780 97.730 98.130 99.890 ;
        RECT 98.610 97.730 98.960 99.890 ;
        RECT 99.440 97.730 99.790 99.890 ;
        RECT 100.270 97.730 100.620 99.890 ;
        RECT 101.100 97.730 101.450 99.890 ;
        RECT 101.930 97.730 102.280 99.890 ;
        RECT 102.760 97.730 103.110 99.890 ;
        RECT 103.590 97.730 103.940 99.890 ;
        RECT 104.420 97.730 104.770 99.890 ;
        RECT 105.250 97.730 105.600 99.890 ;
        RECT 106.080 97.730 106.430 99.890 ;
        RECT 106.910 97.730 107.260 99.890 ;
        RECT 107.740 97.730 108.090 99.890 ;
        RECT 108.570 97.730 108.920 99.890 ;
        RECT 109.400 97.730 109.750 99.890 ;
        RECT 110.230 97.730 110.580 99.890 ;
        RECT 111.060 97.730 111.410 99.890 ;
        RECT 111.890 97.730 112.240 99.890 ;
        RECT 112.720 97.730 113.070 99.890 ;
        RECT 113.550 97.730 113.900 99.890 ;
        RECT 114.380 97.730 114.730 99.890 ;
        RECT 115.210 97.730 115.560 99.890 ;
        RECT 116.040 97.730 116.390 99.890 ;
        RECT 116.870 97.730 117.220 99.890 ;
        RECT 117.700 97.730 118.050 99.890 ;
        RECT 118.530 97.730 118.880 99.890 ;
        RECT 119.360 97.730 119.710 99.890 ;
        RECT 120.190 97.730 120.540 99.890 ;
        RECT 121.020 97.730 121.370 99.890 ;
        RECT 121.850 97.730 122.200 99.890 ;
        RECT 122.680 97.730 123.030 99.890 ;
        RECT 123.510 97.730 123.860 99.890 ;
        RECT 124.340 97.730 124.690 99.890 ;
        RECT 125.170 97.730 125.520 99.890 ;
        RECT 126.000 97.730 126.350 99.890 ;
        RECT 126.830 97.730 127.180 99.890 ;
        RECT 127.660 97.730 128.010 99.890 ;
        RECT 128.490 97.730 128.840 99.890 ;
        RECT 129.320 97.730 129.670 99.890 ;
        RECT 130.150 97.730 130.500 99.890 ;
        RECT 130.980 97.730 131.330 99.890 ;
        RECT 131.810 97.730 132.160 99.890 ;
        RECT 132.640 97.730 132.990 99.890 ;
        RECT 133.470 97.730 133.820 99.890 ;
        RECT 134.300 97.730 134.650 99.890 ;
        RECT 135.130 97.730 135.480 99.890 ;
        RECT 135.960 97.730 136.310 99.890 ;
        RECT 136.790 97.730 137.140 99.890 ;
        RECT 137.620 97.730 137.970 99.890 ;
        RECT 138.450 97.730 138.800 99.890 ;
        RECT 139.280 97.730 139.630 99.890 ;
        RECT 140.110 97.730 140.460 99.890 ;
        RECT 140.940 97.730 141.290 99.890 ;
        RECT 141.770 97.730 142.120 99.890 ;
        RECT 142.600 97.730 142.950 99.890 ;
        RECT 143.430 97.730 143.780 99.890 ;
        RECT 144.260 97.730 144.610 99.890 ;
        RECT 145.090 97.730 145.440 99.890 ;
        RECT 145.920 97.730 146.270 99.890 ;
        RECT 146.750 97.730 147.100 99.890 ;
        RECT 147.580 97.730 147.930 99.890 ;
        RECT 148.410 97.730 148.760 99.890 ;
        RECT 149.240 97.730 149.590 99.890 ;
        RECT 150.070 97.730 150.420 99.890 ;
        RECT 150.900 97.730 151.250 99.890 ;
        RECT 151.730 97.730 152.080 99.890 ;
        RECT 152.560 97.730 152.910 99.890 ;
        RECT 153.390 97.730 153.740 99.890 ;
        RECT 154.220 97.730 154.570 99.890 ;
        RECT 155.050 97.730 155.400 99.890 ;
        RECT 155.880 97.730 156.230 99.890 ;
        RECT 156.710 97.730 157.060 99.890 ;
        RECT 157.540 97.730 157.890 99.890 ;
        RECT 158.370 97.730 158.720 99.890 ;
        RECT 159.200 97.730 159.550 99.890 ;
        RECT 160.030 97.730 160.380 99.890 ;
        RECT 160.860 97.730 161.210 99.890 ;
        RECT 161.690 97.730 162.040 99.890 ;
        RECT 162.520 97.730 162.870 99.890 ;
        RECT 163.350 97.730 163.700 99.890 ;
        RECT 164.180 97.730 164.530 99.890 ;
        RECT 165.010 97.730 165.360 99.890 ;
        RECT 165.840 97.730 166.190 99.890 ;
        RECT 166.670 97.730 167.020 99.890 ;
        RECT 167.500 97.730 167.850 99.890 ;
        RECT 168.330 97.730 168.680 99.890 ;
        RECT 169.160 97.730 169.510 99.890 ;
        RECT 169.990 97.730 170.340 99.890 ;
        RECT 170.820 97.730 171.170 99.890 ;
        RECT 171.650 97.730 172.000 99.890 ;
        RECT 172.480 97.730 172.830 99.890 ;
        RECT 173.310 97.730 173.660 99.890 ;
        RECT 174.140 97.730 174.490 99.890 ;
        RECT 174.970 97.730 175.320 99.890 ;
        RECT 175.800 97.730 176.150 99.890 ;
        RECT 176.630 97.730 176.980 99.890 ;
        RECT 177.460 97.730 177.810 99.890 ;
        RECT 178.290 97.730 178.640 99.890 ;
        RECT 179.120 97.730 179.470 99.890 ;
        RECT 179.950 97.730 180.300 99.890 ;
        RECT 180.780 97.730 181.130 99.890 ;
        RECT 181.610 97.730 181.960 99.890 ;
        RECT 182.440 97.730 182.790 99.890 ;
        RECT 183.270 97.730 183.620 99.890 ;
        RECT 184.100 97.730 184.450 99.890 ;
        RECT 184.930 97.730 185.280 99.890 ;
        RECT 185.760 97.730 186.110 99.890 ;
        RECT 186.590 97.730 186.940 99.890 ;
        RECT 187.420 97.730 187.770 99.890 ;
        RECT 188.250 97.730 188.600 99.890 ;
        RECT 189.080 97.730 189.430 99.890 ;
        RECT 189.910 97.730 190.260 99.890 ;
        RECT 190.740 97.730 191.090 99.890 ;
        RECT 191.570 97.730 191.920 99.890 ;
        RECT 192.400 97.730 192.750 99.890 ;
        RECT 193.230 97.730 193.580 99.890 ;
        RECT 194.060 97.730 194.410 99.890 ;
        RECT 194.890 97.730 195.240 99.890 ;
        RECT 195.720 97.730 196.070 99.890 ;
        RECT 196.550 97.730 196.900 99.890 ;
        RECT 197.380 97.730 197.730 99.890 ;
        RECT 198.210 97.730 198.560 99.890 ;
        RECT 199.040 97.730 199.390 99.890 ;
        RECT 199.870 97.730 200.220 99.890 ;
        RECT 200.700 97.730 201.050 99.890 ;
        RECT 201.530 97.730 201.880 99.890 ;
        RECT 202.360 97.730 202.710 99.890 ;
        RECT 203.190 97.730 203.540 99.890 ;
        RECT 204.020 97.730 204.370 99.890 ;
        RECT 204.850 97.730 205.200 99.890 ;
        RECT 205.680 97.730 206.030 99.890 ;
        RECT 206.510 97.730 206.860 99.890 ;
        RECT 207.340 97.730 207.690 99.890 ;
        RECT 208.170 97.730 208.520 99.890 ;
        RECT 209.000 97.730 209.350 99.890 ;
        RECT 209.830 97.730 210.180 99.890 ;
        RECT 210.660 97.730 211.010 99.890 ;
        RECT 211.490 97.730 211.840 99.890 ;
        RECT 212.320 97.250 212.675 100.500 ;
        RECT 75.275 97.100 212.675 97.250 ;
        RECT 215.625 100.050 228.050 100.500 ;
        RECT 231.045 105.145 271.250 105.495 ;
        RECT 231.045 105.140 249.805 105.145 ;
        RECT 231.045 104.400 231.400 105.140 ;
        RECT 231.670 104.620 232.195 104.945 ;
        RECT 233.495 104.620 234.020 104.945 ;
        RECT 231.800 104.400 231.970 104.415 ;
        RECT 232.280 104.400 232.450 104.415 ;
        RECT 231.045 101.375 232.475 104.400 ;
        RECT 232.760 101.375 232.930 104.415 ;
        RECT 233.240 104.400 233.410 104.415 ;
        RECT 233.720 104.400 233.890 104.415 ;
        RECT 234.290 104.400 236.000 105.140 ;
        RECT 236.270 104.620 236.795 104.945 ;
        RECT 238.095 104.620 238.620 104.945 ;
        RECT 236.400 104.400 236.570 104.415 ;
        RECT 236.880 104.400 237.050 104.415 ;
        RECT 233.225 101.375 237.075 104.400 ;
        RECT 237.360 101.375 237.530 104.415 ;
        RECT 237.840 104.400 238.010 104.415 ;
        RECT 238.320 104.400 238.490 104.415 ;
        RECT 238.890 104.400 240.600 105.140 ;
        RECT 242.570 104.620 242.945 104.945 ;
        RECT 241.000 104.400 241.170 104.415 ;
        RECT 241.480 104.400 241.650 104.415 ;
        RECT 237.825 101.375 241.675 104.400 ;
        RECT 241.960 101.375 242.130 104.415 ;
        RECT 242.440 104.400 242.610 104.415 ;
        RECT 242.920 104.400 243.090 104.415 ;
        RECT 243.490 104.400 245.200 105.140 ;
        RECT 245.470 104.620 245.995 104.945 ;
        RECT 247.295 104.620 247.820 104.945 ;
        RECT 248.090 104.425 249.805 105.140 ;
        RECT 250.080 104.625 250.580 104.950 ;
        RECT 253.830 104.625 254.330 104.950 ;
        RECT 254.605 104.425 271.250 105.145 ;
        RECT 245.600 104.400 245.770 104.415 ;
        RECT 246.080 104.400 246.250 104.415 ;
        RECT 242.425 101.375 246.275 104.400 ;
        RECT 246.560 101.375 246.730 104.415 ;
        RECT 247.040 104.400 247.210 104.415 ;
        RECT 247.520 104.400 247.690 104.415 ;
        RECT 248.090 104.400 250.875 104.425 ;
        RECT 247.025 101.375 250.875 104.400 ;
        RECT 251.160 101.380 251.330 104.420 ;
        RECT 251.640 101.380 251.810 104.420 ;
        RECT 252.120 101.380 252.290 104.420 ;
        RECT 252.600 101.380 252.770 104.420 ;
        RECT 253.080 101.380 253.250 104.420 ;
        RECT 253.525 101.375 271.250 104.425 ;
        RECT 231.045 100.650 231.400 101.375 ;
        RECT 232.445 100.820 233.245 101.195 ;
        RECT 234.290 100.650 236.000 101.375 ;
        RECT 237.045 100.820 237.845 101.195 ;
        RECT 238.890 100.650 240.600 101.375 ;
        RECT 242.095 100.820 242.470 101.195 ;
        RECT 243.490 100.650 245.200 101.375 ;
        RECT 246.245 100.820 247.045 101.195 ;
        RECT 248.090 100.655 249.805 101.375 ;
        RECT 250.830 100.825 253.580 101.200 ;
        RECT 254.605 100.655 271.250 101.375 ;
        RECT 248.090 100.650 271.250 100.655 ;
        RECT 231.045 100.300 271.250 100.650 ;
        RECT 231.045 100.295 234.645 100.300 ;
        RECT 235.645 100.295 239.245 100.300 ;
        RECT 240.245 100.295 243.845 100.300 ;
        RECT 244.845 100.295 248.445 100.300 ;
        RECT 215.625 99.700 254.955 100.050 ;
        RECT 215.625 99.025 231.405 99.700 ;
        RECT 232.450 99.200 233.250 99.525 ;
        RECT 234.295 99.025 236.005 99.700 ;
        RECT 237.050 99.200 237.850 99.525 ;
        RECT 238.895 99.025 240.605 99.700 ;
        RECT 242.100 99.200 242.475 99.525 ;
        RECT 243.495 99.025 245.205 99.700 ;
        RECT 246.250 99.200 247.050 99.525 ;
        RECT 248.095 99.025 249.805 99.700 ;
        RECT 250.830 99.200 253.580 99.525 ;
        RECT 254.605 99.025 254.955 99.700 ;
        RECT 215.625 97.975 232.475 99.025 ;
        RECT 232.765 97.980 232.935 99.020 ;
        RECT 233.225 97.975 237.075 99.025 ;
        RECT 237.365 97.980 237.535 99.020 ;
        RECT 237.825 97.975 241.675 99.025 ;
        RECT 241.965 97.980 242.135 99.020 ;
        RECT 242.425 97.975 246.275 99.025 ;
        RECT 246.565 97.980 246.735 99.020 ;
        RECT 247.025 97.975 250.875 99.025 ;
        RECT 251.160 97.980 251.330 99.020 ;
        RECT 251.640 97.980 251.810 99.020 ;
        RECT 252.120 97.980 252.290 99.020 ;
        RECT 252.600 97.980 252.770 99.020 ;
        RECT 253.080 97.980 253.250 99.020 ;
        RECT 253.525 97.975 254.955 99.025 ;
        RECT 215.625 97.300 231.405 97.975 ;
        RECT 231.675 97.475 232.200 97.800 ;
        RECT 233.500 97.475 234.025 97.800 ;
        RECT 234.295 97.300 236.005 97.975 ;
        RECT 236.275 97.475 236.800 97.800 ;
        RECT 238.100 97.475 238.625 97.800 ;
        RECT 238.895 97.300 240.605 97.975 ;
        RECT 242.575 97.475 242.950 97.800 ;
        RECT 243.495 97.300 245.205 97.975 ;
        RECT 245.475 97.475 246.000 97.800 ;
        RECT 247.300 97.475 247.825 97.800 ;
        RECT 248.095 97.300 249.805 97.975 ;
        RECT 250.080 97.475 250.580 97.800 ;
        RECT 253.830 97.475 254.330 97.800 ;
        RECT 254.605 97.300 254.955 97.975 ;
        RECT 215.625 97.100 254.955 97.300 ;
        RECT 75.275 97.080 212.490 97.100 ;
        RECT 75.275 97.075 97.300 97.080 ;
        RECT 226.800 96.950 254.955 97.100 ;
        RECT 256.625 99.440 271.250 100.300 ;
        RECT 65.075 94.750 70.925 96.325 ;
        RECT 75.280 94.060 226.130 96.395 ;
        RECT 75.280 93.335 76.030 94.060 ;
        RECT 76.260 93.550 77.260 93.720 ;
        RECT 82.710 93.550 83.710 93.720 ;
        RECT 83.930 93.335 86.805 94.060 ;
        RECT 87.010 93.550 88.010 93.720 ;
        RECT 96.040 93.550 97.040 93.720 ;
        RECT 97.255 93.335 100.130 94.060 ;
        RECT 100.335 93.550 101.335 93.720 ;
        RECT 109.365 93.550 110.365 93.720 ;
        RECT 110.580 93.335 113.430 94.060 ;
        RECT 113.660 93.550 114.660 93.720 ;
        RECT 120.110 93.550 121.110 93.720 ;
        RECT 121.330 93.335 124.205 94.060 ;
        RECT 124.410 93.550 125.410 93.720 ;
        RECT 133.440 93.550 134.440 93.720 ;
        RECT 134.655 93.335 137.530 94.060 ;
        RECT 137.735 93.550 138.735 93.720 ;
        RECT 146.765 93.550 147.765 93.720 ;
        RECT 147.980 93.335 150.855 94.060 ;
        RECT 151.060 93.550 152.060 93.720 ;
        RECT 160.090 93.550 161.090 93.720 ;
        RECT 161.305 93.335 164.180 94.060 ;
        RECT 164.385 93.550 165.385 93.720 ;
        RECT 173.415 93.550 174.415 93.720 ;
        RECT 174.630 93.335 177.505 94.060 ;
        RECT 177.710 93.550 178.710 93.720 ;
        RECT 186.740 93.550 187.740 93.720 ;
        RECT 187.955 93.335 190.805 94.060 ;
        RECT 191.035 93.550 192.035 93.720 ;
        RECT 197.485 93.550 198.485 93.720 ;
        RECT 198.705 93.335 201.580 94.060 ;
        RECT 201.785 93.550 202.785 93.720 ;
        RECT 210.815 93.550 211.815 93.720 ;
        RECT 212.030 93.335 214.905 94.060 ;
        RECT 215.110 93.550 216.110 93.720 ;
        RECT 224.140 93.550 225.140 93.720 ;
        RECT 225.355 93.335 226.130 94.060 ;
        RECT 75.280 84.295 76.200 93.335 ;
        RECT 77.320 84.295 77.490 93.335 ;
        RECT 78.610 84.295 78.780 93.335 ;
        RECT 79.900 84.295 80.070 93.335 ;
        RECT 81.190 84.295 81.360 93.335 ;
        RECT 82.480 84.295 82.650 93.335 ;
        RECT 83.770 84.295 86.950 93.335 ;
        RECT 88.070 84.295 88.240 93.335 ;
        RECT 89.360 84.295 89.530 93.335 ;
        RECT 90.650 84.295 90.820 93.335 ;
        RECT 91.940 84.295 92.110 93.335 ;
        RECT 93.230 84.295 93.400 93.335 ;
        RECT 94.520 84.295 94.690 93.335 ;
        RECT 95.810 84.295 95.980 93.335 ;
        RECT 97.100 84.295 100.275 93.335 ;
        RECT 101.395 84.295 101.565 93.335 ;
        RECT 102.685 84.295 102.855 93.335 ;
        RECT 103.975 84.295 104.145 93.335 ;
        RECT 105.265 84.295 105.435 93.335 ;
        RECT 106.555 84.295 106.725 93.335 ;
        RECT 107.845 84.295 108.015 93.335 ;
        RECT 109.135 84.295 109.305 93.335 ;
        RECT 110.425 84.295 113.600 93.335 ;
        RECT 114.720 84.295 114.890 93.335 ;
        RECT 116.010 84.295 116.180 93.335 ;
        RECT 117.300 84.295 117.470 93.335 ;
        RECT 118.590 84.295 118.760 93.335 ;
        RECT 119.880 84.295 120.050 93.335 ;
        RECT 121.170 84.295 124.350 93.335 ;
        RECT 125.470 84.295 125.640 93.335 ;
        RECT 126.760 84.295 126.930 93.335 ;
        RECT 128.050 84.295 128.220 93.335 ;
        RECT 129.340 84.295 129.510 93.335 ;
        RECT 130.630 84.295 130.800 93.335 ;
        RECT 131.920 84.295 132.090 93.335 ;
        RECT 133.210 84.295 133.380 93.335 ;
        RECT 134.500 84.295 137.675 93.335 ;
        RECT 138.795 84.295 138.965 93.335 ;
        RECT 140.085 84.295 140.255 93.335 ;
        RECT 141.375 84.295 141.545 93.335 ;
        RECT 142.665 84.295 142.835 93.335 ;
        RECT 143.955 84.295 144.125 93.335 ;
        RECT 145.245 84.295 145.415 93.335 ;
        RECT 146.535 84.295 146.705 93.335 ;
        RECT 147.825 84.295 151.000 93.335 ;
        RECT 152.120 84.295 152.290 93.335 ;
        RECT 153.410 84.295 153.580 93.335 ;
        RECT 154.700 84.295 154.870 93.335 ;
        RECT 155.990 84.295 156.160 93.335 ;
        RECT 157.280 84.295 157.450 93.335 ;
        RECT 158.570 84.295 158.740 93.335 ;
        RECT 159.860 84.295 160.030 93.335 ;
        RECT 161.150 84.295 164.325 93.335 ;
        RECT 165.445 84.295 165.615 93.335 ;
        RECT 166.735 84.295 166.905 93.335 ;
        RECT 168.025 84.295 168.195 93.335 ;
        RECT 169.315 84.295 169.485 93.335 ;
        RECT 170.605 84.295 170.775 93.335 ;
        RECT 171.895 84.295 172.065 93.335 ;
        RECT 173.185 84.295 173.355 93.335 ;
        RECT 174.475 84.295 177.650 93.335 ;
        RECT 178.770 84.295 178.940 93.335 ;
        RECT 180.060 84.295 180.230 93.335 ;
        RECT 181.350 84.295 181.520 93.335 ;
        RECT 182.640 84.295 182.810 93.335 ;
        RECT 183.930 84.295 184.100 93.335 ;
        RECT 185.220 84.295 185.390 93.335 ;
        RECT 186.510 84.295 186.680 93.335 ;
        RECT 187.800 84.295 190.975 93.335 ;
        RECT 192.095 84.295 192.265 93.335 ;
        RECT 193.385 84.295 193.555 93.335 ;
        RECT 194.675 84.295 194.845 93.335 ;
        RECT 195.965 84.295 196.135 93.335 ;
        RECT 197.255 84.295 197.425 93.335 ;
        RECT 198.545 84.295 201.725 93.335 ;
        RECT 202.845 84.295 203.015 93.335 ;
        RECT 204.135 84.295 204.305 93.335 ;
        RECT 205.425 84.295 205.595 93.335 ;
        RECT 206.715 84.295 206.885 93.335 ;
        RECT 208.005 84.295 208.175 93.335 ;
        RECT 209.295 84.295 209.465 93.335 ;
        RECT 210.585 84.295 210.755 93.335 ;
        RECT 211.875 84.295 215.050 93.335 ;
        RECT 216.170 84.295 216.340 93.335 ;
        RECT 217.460 84.295 217.630 93.335 ;
        RECT 218.750 84.295 218.920 93.335 ;
        RECT 220.040 84.295 220.210 93.335 ;
        RECT 221.330 84.295 221.500 93.335 ;
        RECT 222.620 84.295 222.790 93.335 ;
        RECT 223.910 84.295 224.080 93.335 ;
        RECT 225.200 84.295 226.130 93.335 ;
        RECT 75.280 83.695 76.030 84.295 ;
        RECT 77.550 83.910 78.550 84.080 ;
        RECT 78.840 83.910 79.840 84.080 ;
        RECT 80.130 83.910 81.130 84.080 ;
        RECT 81.420 83.910 82.420 84.080 ;
        RECT 83.930 83.695 86.805 84.295 ;
        RECT 88.300 83.910 89.300 84.080 ;
        RECT 89.590 83.910 90.590 84.080 ;
        RECT 90.880 83.910 91.880 84.080 ;
        RECT 92.170 83.910 93.170 84.080 ;
        RECT 93.460 83.910 94.460 84.080 ;
        RECT 94.750 83.910 95.750 84.080 ;
        RECT 97.255 83.695 100.130 84.295 ;
        RECT 101.625 83.910 102.625 84.080 ;
        RECT 102.915 83.910 103.915 84.080 ;
        RECT 104.205 83.910 105.205 84.080 ;
        RECT 105.495 83.910 106.495 84.080 ;
        RECT 106.785 83.910 107.785 84.080 ;
        RECT 108.075 83.910 109.075 84.080 ;
        RECT 110.580 83.695 113.430 84.295 ;
        RECT 114.950 83.910 115.950 84.080 ;
        RECT 116.240 83.910 117.240 84.080 ;
        RECT 117.530 83.910 118.530 84.080 ;
        RECT 118.820 83.910 119.820 84.080 ;
        RECT 121.330 83.695 124.205 84.295 ;
        RECT 125.700 83.910 126.700 84.080 ;
        RECT 126.990 83.910 127.990 84.080 ;
        RECT 128.280 83.910 129.280 84.080 ;
        RECT 129.570 83.910 130.570 84.080 ;
        RECT 130.860 83.910 131.860 84.080 ;
        RECT 132.150 83.910 133.150 84.080 ;
        RECT 134.655 83.695 137.530 84.295 ;
        RECT 139.025 83.910 140.025 84.080 ;
        RECT 140.315 83.910 141.315 84.080 ;
        RECT 141.605 83.910 142.605 84.080 ;
        RECT 142.895 83.910 143.895 84.080 ;
        RECT 144.185 83.910 145.185 84.080 ;
        RECT 145.475 83.910 146.475 84.080 ;
        RECT 147.980 83.695 150.855 84.295 ;
        RECT 152.350 83.910 153.350 84.080 ;
        RECT 153.640 83.910 154.640 84.080 ;
        RECT 154.930 83.910 155.930 84.080 ;
        RECT 156.220 83.910 157.220 84.080 ;
        RECT 157.510 83.910 158.510 84.080 ;
        RECT 158.800 83.910 159.800 84.080 ;
        RECT 161.305 83.695 164.180 84.295 ;
        RECT 165.675 83.910 166.675 84.080 ;
        RECT 166.965 83.910 167.965 84.080 ;
        RECT 168.255 83.910 169.255 84.080 ;
        RECT 169.545 83.910 170.545 84.080 ;
        RECT 170.835 83.910 171.835 84.080 ;
        RECT 172.125 83.910 173.125 84.080 ;
        RECT 174.630 83.695 177.505 84.295 ;
        RECT 179.000 83.910 180.000 84.080 ;
        RECT 180.290 83.910 181.290 84.080 ;
        RECT 181.580 83.910 182.580 84.080 ;
        RECT 182.870 83.910 183.870 84.080 ;
        RECT 184.160 83.910 185.160 84.080 ;
        RECT 185.450 83.910 186.450 84.080 ;
        RECT 187.955 83.695 190.805 84.295 ;
        RECT 192.325 83.910 193.325 84.080 ;
        RECT 193.615 83.910 194.615 84.080 ;
        RECT 194.905 83.910 195.905 84.080 ;
        RECT 196.195 83.910 197.195 84.080 ;
        RECT 198.705 83.695 201.580 84.295 ;
        RECT 203.075 83.910 204.075 84.080 ;
        RECT 204.365 83.910 205.365 84.080 ;
        RECT 205.655 83.910 206.655 84.080 ;
        RECT 206.945 83.910 207.945 84.080 ;
        RECT 208.235 83.910 209.235 84.080 ;
        RECT 209.525 83.910 210.525 84.080 ;
        RECT 212.030 83.695 214.905 84.295 ;
        RECT 216.400 83.910 217.400 84.080 ;
        RECT 217.690 83.910 218.690 84.080 ;
        RECT 218.980 83.910 219.980 84.080 ;
        RECT 220.270 83.910 221.270 84.080 ;
        RECT 221.560 83.910 222.560 84.080 ;
        RECT 222.850 83.910 223.850 84.080 ;
        RECT 225.355 83.695 226.130 84.295 ;
        RECT 72.725 82.575 73.450 83.675 ;
        RECT 75.280 83.400 226.130 83.695 ;
        RECT 75.280 83.395 76.030 83.400 ;
        RECT 83.930 83.395 86.805 83.400 ;
        RECT 97.255 83.395 100.130 83.400 ;
        RECT 110.580 83.395 113.430 83.400 ;
        RECT 121.330 83.395 124.205 83.400 ;
        RECT 134.655 83.395 137.530 83.400 ;
        RECT 147.980 83.395 150.855 83.400 ;
        RECT 161.305 83.395 164.180 83.400 ;
        RECT 174.630 83.395 177.505 83.400 ;
        RECT 187.955 83.395 190.805 83.400 ;
        RECT 198.705 83.395 201.580 83.400 ;
        RECT 212.030 83.395 214.905 83.400 ;
        RECT 225.355 83.395 226.130 83.400 ;
        RECT 226.800 90.750 228.050 96.950 ;
        RECT 231.050 96.200 233.700 96.205 ;
        RECT 231.050 95.850 254.955 96.200 ;
        RECT 231.050 91.360 231.425 95.850 ;
        RECT 233.325 95.845 254.955 95.850 ;
        RECT 233.325 95.840 249.805 95.845 ;
        RECT 231.950 95.305 232.800 95.680 ;
        RECT 231.810 92.085 231.980 95.125 ;
        RECT 232.290 92.085 232.460 95.125 ;
        RECT 232.770 92.085 232.940 95.125 ;
        RECT 233.325 95.100 236.000 95.840 ;
        RECT 236.270 95.320 236.795 95.645 ;
        RECT 238.095 95.320 238.620 95.645 ;
        RECT 236.400 95.100 236.570 95.115 ;
        RECT 236.880 95.100 237.050 95.115 ;
        RECT 233.325 92.075 237.075 95.100 ;
        RECT 237.360 92.075 237.530 95.115 ;
        RECT 237.840 95.100 238.010 95.115 ;
        RECT 238.320 95.100 238.490 95.115 ;
        RECT 238.890 95.100 240.600 95.840 ;
        RECT 242.570 95.320 242.945 95.645 ;
        RECT 241.000 95.100 241.170 95.115 ;
        RECT 241.480 95.100 241.650 95.115 ;
        RECT 237.825 92.075 241.675 95.100 ;
        RECT 241.960 92.075 242.130 95.115 ;
        RECT 242.440 95.100 242.610 95.115 ;
        RECT 242.920 95.100 243.090 95.115 ;
        RECT 243.490 95.100 245.200 95.840 ;
        RECT 245.470 95.320 245.995 95.645 ;
        RECT 247.295 95.320 247.820 95.645 ;
        RECT 248.090 95.125 249.805 95.840 ;
        RECT 250.080 95.325 250.580 95.650 ;
        RECT 253.830 95.325 254.330 95.650 ;
        RECT 254.605 95.125 254.955 95.845 ;
        RECT 245.600 95.100 245.770 95.115 ;
        RECT 246.080 95.100 246.250 95.115 ;
        RECT 242.425 92.075 246.275 95.100 ;
        RECT 246.560 92.075 246.730 95.115 ;
        RECT 247.040 95.100 247.210 95.115 ;
        RECT 247.520 95.100 247.690 95.115 ;
        RECT 248.090 95.100 250.875 95.125 ;
        RECT 247.025 92.075 250.875 95.100 ;
        RECT 251.160 92.080 251.330 95.120 ;
        RECT 251.640 92.080 251.810 95.120 ;
        RECT 252.120 92.080 252.290 95.120 ;
        RECT 252.600 92.080 252.770 95.120 ;
        RECT 253.080 92.080 253.250 95.120 ;
        RECT 253.525 92.075 254.955 95.125 ;
        RECT 256.625 94.950 256.975 99.440 ;
        RECT 257.540 98.895 259.290 99.270 ;
        RECT 268.590 98.895 270.340 99.270 ;
        RECT 257.375 95.675 257.545 98.715 ;
        RECT 257.855 95.675 258.025 98.715 ;
        RECT 258.335 95.675 258.505 98.715 ;
        RECT 258.815 95.675 258.985 98.715 ;
        RECT 259.295 95.675 259.465 98.715 ;
        RECT 259.775 95.675 259.945 98.715 ;
        RECT 260.255 95.675 260.425 98.715 ;
        RECT 260.735 95.675 260.905 98.715 ;
        RECT 261.215 95.675 261.385 98.715 ;
        RECT 261.695 95.675 261.865 98.715 ;
        RECT 262.175 95.675 262.345 98.715 ;
        RECT 262.655 95.675 262.825 98.715 ;
        RECT 263.135 95.675 263.305 98.715 ;
        RECT 263.615 95.675 263.785 98.715 ;
        RECT 264.095 95.675 264.265 98.715 ;
        RECT 264.575 95.675 264.745 98.715 ;
        RECT 265.055 95.675 265.225 98.715 ;
        RECT 265.535 95.675 265.705 98.715 ;
        RECT 266.015 95.675 266.185 98.715 ;
        RECT 266.495 95.675 266.665 98.715 ;
        RECT 266.975 95.675 267.145 98.715 ;
        RECT 267.455 95.675 267.625 98.715 ;
        RECT 267.935 95.675 268.105 98.715 ;
        RECT 268.415 95.675 268.585 98.715 ;
        RECT 268.895 95.675 269.065 98.715 ;
        RECT 269.375 95.675 269.545 98.715 ;
        RECT 269.855 95.675 270.025 98.715 ;
        RECT 270.335 95.675 270.505 98.715 ;
        RECT 259.465 95.120 268.415 95.495 ;
        RECT 270.900 94.950 271.250 99.440 ;
        RECT 256.625 94.600 271.250 94.950 ;
        RECT 233.325 91.360 236.000 92.075 ;
        RECT 237.045 91.520 237.845 91.895 ;
        RECT 231.050 91.350 236.000 91.360 ;
        RECT 238.890 91.350 240.600 92.075 ;
        RECT 242.095 91.520 242.470 91.895 ;
        RECT 243.490 91.350 245.200 92.075 ;
        RECT 246.245 91.520 247.045 91.895 ;
        RECT 248.090 91.355 249.805 92.075 ;
        RECT 250.830 91.525 253.580 91.900 ;
        RECT 254.605 91.355 254.955 92.075 ;
        RECT 248.090 91.350 254.955 91.355 ;
        RECT 231.050 91.005 254.955 91.350 ;
        RECT 233.325 91.000 254.955 91.005 ;
        RECT 256.625 94.000 271.250 94.350 ;
        RECT 256.625 91.600 256.975 94.000 ;
        RECT 257.540 93.500 259.290 93.825 ;
        RECT 268.590 93.500 270.340 93.825 ;
        RECT 257.375 92.280 257.545 93.320 ;
        RECT 257.855 92.280 258.025 93.320 ;
        RECT 258.335 92.280 258.505 93.320 ;
        RECT 258.815 92.280 258.985 93.320 ;
        RECT 259.295 92.280 259.465 93.320 ;
        RECT 259.775 92.280 259.945 93.320 ;
        RECT 260.255 92.280 260.425 93.320 ;
        RECT 260.735 92.280 260.905 93.320 ;
        RECT 261.215 92.280 261.385 93.320 ;
        RECT 261.695 92.280 261.865 93.320 ;
        RECT 262.175 92.280 262.345 93.320 ;
        RECT 262.655 92.280 262.825 93.320 ;
        RECT 263.135 92.280 263.305 93.320 ;
        RECT 263.615 92.280 263.785 93.320 ;
        RECT 264.095 92.280 264.265 93.320 ;
        RECT 264.575 92.280 264.745 93.320 ;
        RECT 265.055 92.280 265.225 93.320 ;
        RECT 265.535 92.280 265.705 93.320 ;
        RECT 266.015 92.280 266.185 93.320 ;
        RECT 266.495 92.280 266.665 93.320 ;
        RECT 266.975 92.280 267.145 93.320 ;
        RECT 267.455 92.280 267.625 93.320 ;
        RECT 267.935 92.280 268.105 93.320 ;
        RECT 268.415 92.280 268.585 93.320 ;
        RECT 268.895 92.280 269.065 93.320 ;
        RECT 269.375 92.280 269.545 93.320 ;
        RECT 269.855 92.280 270.025 93.320 ;
        RECT 270.335 92.280 270.505 93.320 ;
        RECT 259.465 91.775 268.415 92.100 ;
        RECT 270.900 91.600 271.250 94.000 ;
        RECT 235.645 90.995 239.245 91.000 ;
        RECT 240.245 90.995 243.845 91.000 ;
        RECT 244.845 90.995 248.445 91.000 ;
        RECT 256.625 90.750 271.250 91.600 ;
        RECT 226.800 90.400 271.250 90.750 ;
        RECT 226.800 88.000 231.425 90.400 ;
        RECT 233.325 89.725 236.005 90.400 ;
        RECT 237.050 89.900 237.850 90.225 ;
        RECT 238.895 89.725 240.605 90.400 ;
        RECT 242.100 89.900 242.475 90.225 ;
        RECT 243.495 89.725 245.205 90.400 ;
        RECT 246.250 89.900 247.050 90.225 ;
        RECT 248.095 89.725 249.805 90.400 ;
        RECT 250.830 89.900 253.580 90.225 ;
        RECT 254.605 89.725 271.250 90.400 ;
        RECT 231.810 88.680 231.980 89.720 ;
        RECT 232.290 88.680 232.460 89.720 ;
        RECT 232.770 88.680 232.940 89.720 ;
        RECT 233.325 88.675 237.075 89.725 ;
        RECT 237.365 88.680 237.535 89.720 ;
        RECT 237.825 88.675 241.675 89.725 ;
        RECT 241.965 88.680 242.135 89.720 ;
        RECT 242.425 88.675 246.275 89.725 ;
        RECT 246.565 88.680 246.735 89.720 ;
        RECT 247.025 88.675 250.875 89.725 ;
        RECT 251.160 88.680 251.330 89.720 ;
        RECT 251.640 88.680 251.810 89.720 ;
        RECT 252.120 88.680 252.290 89.720 ;
        RECT 252.600 88.680 252.770 89.720 ;
        RECT 253.080 88.680 253.250 89.720 ;
        RECT 253.525 88.675 271.250 89.725 ;
        RECT 231.950 88.175 232.800 88.500 ;
        RECT 233.325 88.000 236.005 88.675 ;
        RECT 236.275 88.175 236.800 88.500 ;
        RECT 238.100 88.175 238.625 88.500 ;
        RECT 238.895 88.000 240.605 88.675 ;
        RECT 242.575 88.175 242.950 88.500 ;
        RECT 243.495 88.000 245.205 88.675 ;
        RECT 245.475 88.175 246.000 88.500 ;
        RECT 247.300 88.175 247.825 88.500 ;
        RECT 248.095 88.000 249.805 88.675 ;
        RECT 250.080 88.175 250.580 88.500 ;
        RECT 253.830 88.175 254.330 88.500 ;
        RECT 254.605 88.000 271.250 88.675 ;
        RECT 226.800 86.800 271.250 88.000 ;
        RECT 75.280 82.545 226.130 82.845 ;
        RECT 75.280 81.990 76.030 82.545 ;
        RECT 77.550 82.160 78.550 82.330 ;
        RECT 78.840 82.160 79.840 82.330 ;
        RECT 80.130 82.160 81.130 82.330 ;
        RECT 81.420 82.160 82.420 82.330 ;
        RECT 83.930 81.990 86.805 82.545 ;
        RECT 88.300 82.160 89.300 82.330 ;
        RECT 89.590 82.160 90.590 82.330 ;
        RECT 90.880 82.160 91.880 82.330 ;
        RECT 92.170 82.160 93.170 82.330 ;
        RECT 93.460 82.160 94.460 82.330 ;
        RECT 94.750 82.160 95.750 82.330 ;
        RECT 97.255 81.990 100.130 82.545 ;
        RECT 101.625 82.160 102.625 82.330 ;
        RECT 102.915 82.160 103.915 82.330 ;
        RECT 104.205 82.160 105.205 82.330 ;
        RECT 105.495 82.160 106.495 82.330 ;
        RECT 106.785 82.160 107.785 82.330 ;
        RECT 108.075 82.160 109.075 82.330 ;
        RECT 110.580 81.990 113.430 82.545 ;
        RECT 114.950 82.160 115.950 82.330 ;
        RECT 116.240 82.160 117.240 82.330 ;
        RECT 117.530 82.160 118.530 82.330 ;
        RECT 118.820 82.160 119.820 82.330 ;
        RECT 121.330 81.990 124.205 82.545 ;
        RECT 125.700 82.160 126.700 82.330 ;
        RECT 126.990 82.160 127.990 82.330 ;
        RECT 128.280 82.160 129.280 82.330 ;
        RECT 129.570 82.160 130.570 82.330 ;
        RECT 130.860 82.160 131.860 82.330 ;
        RECT 132.150 82.160 133.150 82.330 ;
        RECT 134.655 81.990 137.530 82.545 ;
        RECT 139.025 82.160 140.025 82.330 ;
        RECT 140.315 82.160 141.315 82.330 ;
        RECT 141.605 82.160 142.605 82.330 ;
        RECT 142.895 82.160 143.895 82.330 ;
        RECT 144.185 82.160 145.185 82.330 ;
        RECT 145.475 82.160 146.475 82.330 ;
        RECT 147.980 81.990 150.855 82.545 ;
        RECT 152.350 82.160 153.350 82.330 ;
        RECT 153.640 82.160 154.640 82.330 ;
        RECT 154.930 82.160 155.930 82.330 ;
        RECT 156.220 82.160 157.220 82.330 ;
        RECT 157.510 82.160 158.510 82.330 ;
        RECT 158.800 82.160 159.800 82.330 ;
        RECT 161.305 81.990 164.180 82.545 ;
        RECT 165.675 82.160 166.675 82.330 ;
        RECT 166.965 82.160 167.965 82.330 ;
        RECT 168.255 82.160 169.255 82.330 ;
        RECT 169.545 82.160 170.545 82.330 ;
        RECT 170.835 82.160 171.835 82.330 ;
        RECT 172.125 82.160 173.125 82.330 ;
        RECT 174.630 81.990 177.505 82.545 ;
        RECT 179.000 82.160 180.000 82.330 ;
        RECT 180.290 82.160 181.290 82.330 ;
        RECT 181.580 82.160 182.580 82.330 ;
        RECT 182.870 82.160 183.870 82.330 ;
        RECT 184.160 82.160 185.160 82.330 ;
        RECT 185.450 82.160 186.450 82.330 ;
        RECT 187.955 81.990 190.805 82.545 ;
        RECT 192.325 82.160 193.325 82.330 ;
        RECT 193.615 82.160 194.615 82.330 ;
        RECT 194.905 82.160 195.905 82.330 ;
        RECT 196.195 82.160 197.195 82.330 ;
        RECT 198.705 81.990 201.580 82.545 ;
        RECT 203.075 82.160 204.075 82.330 ;
        RECT 204.365 82.160 205.365 82.330 ;
        RECT 205.655 82.160 206.655 82.330 ;
        RECT 206.945 82.160 207.945 82.330 ;
        RECT 208.235 82.160 209.235 82.330 ;
        RECT 209.525 82.160 210.525 82.330 ;
        RECT 212.030 81.990 214.905 82.545 ;
        RECT 216.400 82.160 217.400 82.330 ;
        RECT 217.690 82.160 218.690 82.330 ;
        RECT 218.980 82.160 219.980 82.330 ;
        RECT 220.270 82.160 221.270 82.330 ;
        RECT 221.560 82.160 222.560 82.330 ;
        RECT 222.850 82.160 223.850 82.330 ;
        RECT 225.355 82.000 226.130 82.545 ;
        RECT 226.800 82.000 228.050 86.800 ;
        RECT 231.050 84.645 271.250 85.500 ;
        RECT 225.355 81.990 228.050 82.000 ;
        RECT 75.280 78.950 76.200 81.990 ;
        RECT 77.320 78.950 77.490 81.990 ;
        RECT 78.610 78.950 78.780 81.990 ;
        RECT 79.900 78.950 80.070 81.990 ;
        RECT 81.190 78.950 81.360 81.990 ;
        RECT 82.480 78.950 82.650 81.990 ;
        RECT 83.770 78.950 86.950 81.990 ;
        RECT 88.070 78.950 88.240 81.990 ;
        RECT 89.360 78.950 89.530 81.990 ;
        RECT 90.650 78.950 90.820 81.990 ;
        RECT 91.940 78.950 92.110 81.990 ;
        RECT 93.230 78.950 93.400 81.990 ;
        RECT 94.520 78.950 94.690 81.990 ;
        RECT 95.810 78.950 95.980 81.990 ;
        RECT 97.100 78.950 100.275 81.990 ;
        RECT 101.395 78.950 101.565 81.990 ;
        RECT 102.685 78.950 102.855 81.990 ;
        RECT 103.975 78.950 104.145 81.990 ;
        RECT 105.265 78.950 105.435 81.990 ;
        RECT 106.555 78.950 106.725 81.990 ;
        RECT 107.845 78.950 108.015 81.990 ;
        RECT 109.135 78.950 109.305 81.990 ;
        RECT 110.425 78.950 113.600 81.990 ;
        RECT 114.720 78.950 114.890 81.990 ;
        RECT 116.010 78.950 116.180 81.990 ;
        RECT 117.300 78.950 117.470 81.990 ;
        RECT 118.590 78.950 118.760 81.990 ;
        RECT 119.880 78.950 120.050 81.990 ;
        RECT 121.170 78.950 124.350 81.990 ;
        RECT 125.470 78.950 125.640 81.990 ;
        RECT 126.760 78.950 126.930 81.990 ;
        RECT 128.050 78.950 128.220 81.990 ;
        RECT 129.340 78.950 129.510 81.990 ;
        RECT 130.630 78.950 130.800 81.990 ;
        RECT 131.920 78.950 132.090 81.990 ;
        RECT 133.210 78.950 133.380 81.990 ;
        RECT 134.500 78.950 137.675 81.990 ;
        RECT 138.795 78.950 138.965 81.990 ;
        RECT 140.085 78.950 140.255 81.990 ;
        RECT 141.375 78.950 141.545 81.990 ;
        RECT 142.665 78.950 142.835 81.990 ;
        RECT 143.955 78.950 144.125 81.990 ;
        RECT 145.245 78.950 145.415 81.990 ;
        RECT 146.535 78.950 146.705 81.990 ;
        RECT 147.825 78.950 151.000 81.990 ;
        RECT 152.120 78.950 152.290 81.990 ;
        RECT 153.410 78.950 153.580 81.990 ;
        RECT 154.700 78.950 154.870 81.990 ;
        RECT 155.990 78.950 156.160 81.990 ;
        RECT 157.280 78.950 157.450 81.990 ;
        RECT 158.570 78.950 158.740 81.990 ;
        RECT 159.860 78.950 160.030 81.990 ;
        RECT 161.150 78.950 164.325 81.990 ;
        RECT 165.445 78.950 165.615 81.990 ;
        RECT 166.735 78.950 166.905 81.990 ;
        RECT 168.025 78.950 168.195 81.990 ;
        RECT 169.315 78.950 169.485 81.990 ;
        RECT 170.605 78.950 170.775 81.990 ;
        RECT 171.895 78.950 172.065 81.990 ;
        RECT 173.185 78.950 173.355 81.990 ;
        RECT 174.475 78.950 177.650 81.990 ;
        RECT 178.770 78.950 178.940 81.990 ;
        RECT 180.060 78.950 180.230 81.990 ;
        RECT 181.350 78.950 181.520 81.990 ;
        RECT 182.640 78.950 182.810 81.990 ;
        RECT 183.930 78.950 184.100 81.990 ;
        RECT 185.220 78.950 185.390 81.990 ;
        RECT 186.510 78.950 186.680 81.990 ;
        RECT 187.800 78.950 190.975 81.990 ;
        RECT 192.095 78.950 192.265 81.990 ;
        RECT 193.385 78.950 193.555 81.990 ;
        RECT 194.675 78.950 194.845 81.990 ;
        RECT 195.965 78.950 196.135 81.990 ;
        RECT 197.255 78.950 197.425 81.990 ;
        RECT 198.545 78.950 201.725 81.990 ;
        RECT 202.845 78.950 203.015 81.990 ;
        RECT 204.135 78.950 204.305 81.990 ;
        RECT 205.425 78.950 205.595 81.990 ;
        RECT 206.715 78.950 206.885 81.990 ;
        RECT 208.005 78.950 208.175 81.990 ;
        RECT 209.295 78.950 209.465 81.990 ;
        RECT 210.585 78.950 210.755 81.990 ;
        RECT 211.875 78.950 215.050 81.990 ;
        RECT 216.170 78.950 216.340 81.990 ;
        RECT 217.460 78.950 217.630 81.990 ;
        RECT 218.750 78.950 218.920 81.990 ;
        RECT 220.040 78.950 220.210 81.990 ;
        RECT 221.330 78.950 221.500 81.990 ;
        RECT 222.620 78.950 222.790 81.990 ;
        RECT 223.910 78.950 224.080 81.990 ;
        RECT 225.200 79.200 228.050 81.990 ;
        RECT 231.045 84.295 271.250 84.645 ;
        RECT 231.045 84.290 249.805 84.295 ;
        RECT 231.045 83.550 231.400 84.290 ;
        RECT 231.670 83.770 232.195 84.095 ;
        RECT 233.495 83.770 234.020 84.095 ;
        RECT 231.800 83.550 231.970 83.565 ;
        RECT 232.280 83.550 232.450 83.565 ;
        RECT 231.045 80.525 232.475 83.550 ;
        RECT 232.760 80.525 232.930 83.565 ;
        RECT 233.240 83.550 233.410 83.565 ;
        RECT 233.720 83.550 233.890 83.565 ;
        RECT 234.290 83.550 236.000 84.290 ;
        RECT 236.270 83.770 236.795 84.095 ;
        RECT 238.095 83.770 238.620 84.095 ;
        RECT 236.400 83.550 236.570 83.565 ;
        RECT 236.880 83.550 237.050 83.565 ;
        RECT 233.225 80.525 237.075 83.550 ;
        RECT 237.360 80.525 237.530 83.565 ;
        RECT 237.840 83.550 238.010 83.565 ;
        RECT 238.320 83.550 238.490 83.565 ;
        RECT 238.890 83.550 240.600 84.290 ;
        RECT 242.570 83.770 242.945 84.095 ;
        RECT 241.000 83.550 241.170 83.565 ;
        RECT 241.480 83.550 241.650 83.565 ;
        RECT 237.825 80.525 241.675 83.550 ;
        RECT 241.960 80.525 242.130 83.565 ;
        RECT 242.440 83.550 242.610 83.565 ;
        RECT 242.920 83.550 243.090 83.565 ;
        RECT 243.490 83.550 245.200 84.290 ;
        RECT 245.470 83.770 245.995 84.095 ;
        RECT 247.295 83.770 247.820 84.095 ;
        RECT 248.090 83.575 249.805 84.290 ;
        RECT 250.080 83.775 250.580 84.100 ;
        RECT 253.830 83.775 254.330 84.100 ;
        RECT 254.605 83.575 271.250 84.295 ;
        RECT 245.600 83.550 245.770 83.565 ;
        RECT 246.080 83.550 246.250 83.565 ;
        RECT 242.425 80.525 246.275 83.550 ;
        RECT 246.560 80.525 246.730 83.565 ;
        RECT 247.040 83.550 247.210 83.565 ;
        RECT 247.520 83.550 247.690 83.565 ;
        RECT 248.090 83.550 250.875 83.575 ;
        RECT 247.025 80.525 250.875 83.550 ;
        RECT 251.160 80.530 251.330 83.570 ;
        RECT 251.640 80.530 251.810 83.570 ;
        RECT 252.120 80.530 252.290 83.570 ;
        RECT 252.600 80.530 252.770 83.570 ;
        RECT 253.080 80.530 253.250 83.570 ;
        RECT 253.525 80.525 271.250 83.575 ;
        RECT 231.045 79.800 231.400 80.525 ;
        RECT 232.445 79.970 233.245 80.345 ;
        RECT 234.290 79.800 236.000 80.525 ;
        RECT 237.045 79.970 237.845 80.345 ;
        RECT 238.890 79.800 240.600 80.525 ;
        RECT 242.095 79.970 242.470 80.345 ;
        RECT 243.490 79.800 245.200 80.525 ;
        RECT 246.245 79.970 247.045 80.345 ;
        RECT 248.090 79.805 249.805 80.525 ;
        RECT 250.830 79.975 253.580 80.350 ;
        RECT 254.605 79.805 271.250 80.525 ;
        RECT 248.090 79.800 271.250 79.805 ;
        RECT 231.045 79.450 271.250 79.800 ;
        RECT 231.045 79.445 234.645 79.450 ;
        RECT 235.645 79.445 239.245 79.450 ;
        RECT 240.245 79.445 243.845 79.450 ;
        RECT 244.845 79.445 248.445 79.450 ;
        RECT 225.200 78.950 254.955 79.200 ;
        RECT 75.280 78.270 76.030 78.950 ;
        RECT 76.260 78.610 77.260 78.780 ;
        RECT 82.710 78.610 83.710 78.780 ;
        RECT 83.930 78.270 86.805 78.950 ;
        RECT 87.010 78.610 88.010 78.780 ;
        RECT 96.040 78.610 97.040 78.780 ;
        RECT 97.255 78.270 100.130 78.950 ;
        RECT 100.335 78.610 101.335 78.780 ;
        RECT 109.365 78.610 110.365 78.780 ;
        RECT 110.580 78.270 113.430 78.950 ;
        RECT 113.660 78.610 114.660 78.780 ;
        RECT 120.110 78.610 121.110 78.780 ;
        RECT 121.330 78.270 124.205 78.950 ;
        RECT 124.410 78.610 125.410 78.780 ;
        RECT 133.440 78.610 134.440 78.780 ;
        RECT 134.655 78.270 137.530 78.950 ;
        RECT 137.735 78.610 138.735 78.780 ;
        RECT 146.765 78.610 147.765 78.780 ;
        RECT 147.980 78.270 150.855 78.950 ;
        RECT 151.060 78.610 152.060 78.780 ;
        RECT 160.090 78.610 161.090 78.780 ;
        RECT 161.305 78.270 164.180 78.950 ;
        RECT 164.385 78.610 165.385 78.780 ;
        RECT 173.415 78.610 174.415 78.780 ;
        RECT 174.630 78.270 177.505 78.950 ;
        RECT 177.710 78.610 178.710 78.780 ;
        RECT 186.740 78.610 187.740 78.780 ;
        RECT 187.955 78.270 190.805 78.950 ;
        RECT 191.035 78.610 192.035 78.780 ;
        RECT 197.485 78.610 198.485 78.780 ;
        RECT 198.705 78.270 201.580 78.950 ;
        RECT 201.785 78.610 202.785 78.780 ;
        RECT 210.815 78.610 211.815 78.780 ;
        RECT 212.030 78.270 214.905 78.950 ;
        RECT 225.355 78.850 254.955 78.950 ;
        RECT 215.110 78.610 216.110 78.780 ;
        RECT 224.140 78.610 225.140 78.780 ;
        RECT 225.355 78.270 231.405 78.850 ;
        RECT 232.450 78.350 233.250 78.675 ;
        RECT 75.280 78.175 231.405 78.270 ;
        RECT 234.295 78.175 236.005 78.850 ;
        RECT 237.050 78.350 237.850 78.675 ;
        RECT 238.895 78.175 240.605 78.850 ;
        RECT 242.100 78.350 242.475 78.675 ;
        RECT 243.495 78.175 245.205 78.850 ;
        RECT 246.250 78.350 247.050 78.675 ;
        RECT 248.095 78.175 249.805 78.850 ;
        RECT 250.830 78.350 253.580 78.675 ;
        RECT 254.605 78.175 254.955 78.850 ;
        RECT 75.280 77.125 232.475 78.175 ;
        RECT 232.765 77.130 232.935 78.170 ;
        RECT 233.225 77.125 237.075 78.175 ;
        RECT 237.365 77.130 237.535 78.170 ;
        RECT 237.825 77.125 241.675 78.175 ;
        RECT 241.965 77.130 242.135 78.170 ;
        RECT 242.425 77.125 246.275 78.175 ;
        RECT 246.565 77.130 246.735 78.170 ;
        RECT 247.025 77.125 250.875 78.175 ;
        RECT 251.160 77.130 251.330 78.170 ;
        RECT 251.640 77.130 251.810 78.170 ;
        RECT 252.120 77.130 252.290 78.170 ;
        RECT 252.600 77.130 252.770 78.170 ;
        RECT 253.080 77.130 253.250 78.170 ;
        RECT 253.525 77.125 254.955 78.175 ;
        RECT 75.280 76.450 231.405 77.125 ;
        RECT 231.675 76.625 232.200 76.950 ;
        RECT 233.500 76.625 234.025 76.950 ;
        RECT 234.295 76.450 236.005 77.125 ;
        RECT 236.275 76.625 236.800 76.950 ;
        RECT 238.100 76.625 238.625 76.950 ;
        RECT 238.895 76.450 240.605 77.125 ;
        RECT 242.575 76.625 242.950 76.950 ;
        RECT 243.495 76.450 245.205 77.125 ;
        RECT 245.475 76.625 246.000 76.950 ;
        RECT 247.300 76.625 247.825 76.950 ;
        RECT 248.095 76.450 249.805 77.125 ;
        RECT 250.080 76.625 250.580 76.950 ;
        RECT 253.830 76.625 254.330 76.950 ;
        RECT 254.605 76.450 254.955 77.125 ;
        RECT 75.280 76.100 254.955 76.450 ;
        RECT 256.625 78.590 271.250 79.450 ;
        RECT 75.280 75.945 228.050 76.100 ;
        RECT 97.130 75.300 212.490 75.315 ;
        RECT 75.275 75.145 212.675 75.300 ;
        RECT 75.275 68.025 97.300 75.145 ;
        RECT 97.780 72.505 98.130 74.665 ;
        RECT 98.610 72.505 98.960 74.665 ;
        RECT 99.440 72.505 99.790 74.665 ;
        RECT 100.270 72.505 100.620 74.665 ;
        RECT 101.100 72.505 101.450 74.665 ;
        RECT 101.930 72.505 102.280 74.665 ;
        RECT 102.760 72.505 103.110 74.665 ;
        RECT 103.590 72.505 103.940 74.665 ;
        RECT 104.420 72.505 104.770 74.665 ;
        RECT 105.250 72.505 105.600 74.665 ;
        RECT 106.080 72.505 106.430 74.665 ;
        RECT 106.910 72.505 107.260 74.665 ;
        RECT 107.740 72.505 108.090 74.665 ;
        RECT 108.570 72.505 108.920 74.665 ;
        RECT 109.400 72.505 109.750 74.665 ;
        RECT 110.230 72.505 110.580 74.665 ;
        RECT 111.060 72.505 111.410 74.665 ;
        RECT 111.890 72.505 112.240 74.665 ;
        RECT 112.720 72.505 113.070 74.665 ;
        RECT 113.550 72.505 113.900 74.665 ;
        RECT 114.380 72.505 114.730 74.665 ;
        RECT 115.210 72.505 115.560 74.665 ;
        RECT 116.040 72.505 116.390 74.665 ;
        RECT 116.870 72.505 117.220 74.665 ;
        RECT 117.700 72.505 118.050 74.665 ;
        RECT 118.530 72.505 118.880 74.665 ;
        RECT 119.360 72.505 119.710 74.665 ;
        RECT 120.190 72.505 120.540 74.665 ;
        RECT 121.020 72.505 121.370 74.665 ;
        RECT 121.850 72.505 122.200 74.665 ;
        RECT 122.680 72.505 123.030 74.665 ;
        RECT 123.510 72.505 123.860 74.665 ;
        RECT 124.340 72.505 124.690 74.665 ;
        RECT 125.170 72.505 125.520 74.665 ;
        RECT 126.000 72.505 126.350 74.665 ;
        RECT 126.830 72.505 127.180 74.665 ;
        RECT 127.660 72.505 128.010 74.665 ;
        RECT 128.490 72.505 128.840 74.665 ;
        RECT 129.320 72.505 129.670 74.665 ;
        RECT 130.150 72.505 130.500 74.665 ;
        RECT 130.980 72.505 131.330 74.665 ;
        RECT 131.810 72.505 132.160 74.665 ;
        RECT 132.640 72.505 132.990 74.665 ;
        RECT 133.470 72.505 133.820 74.665 ;
        RECT 134.300 72.505 134.650 74.665 ;
        RECT 135.130 72.505 135.480 74.665 ;
        RECT 135.960 72.505 136.310 74.665 ;
        RECT 136.790 72.505 137.140 74.665 ;
        RECT 137.620 72.505 137.970 74.665 ;
        RECT 138.450 72.505 138.800 74.665 ;
        RECT 139.280 72.505 139.630 74.665 ;
        RECT 140.110 72.505 140.460 74.665 ;
        RECT 140.940 72.505 141.290 74.665 ;
        RECT 141.770 72.505 142.120 74.665 ;
        RECT 142.600 72.505 142.950 74.665 ;
        RECT 143.430 72.505 143.780 74.665 ;
        RECT 144.260 72.505 144.610 74.665 ;
        RECT 145.090 72.505 145.440 74.665 ;
        RECT 145.920 72.505 146.270 74.665 ;
        RECT 146.750 72.505 147.100 74.665 ;
        RECT 147.580 72.505 147.930 74.665 ;
        RECT 148.410 72.505 148.760 74.665 ;
        RECT 149.240 72.505 149.590 74.665 ;
        RECT 150.070 72.505 150.420 74.665 ;
        RECT 150.900 72.505 151.250 74.665 ;
        RECT 151.730 72.505 152.080 74.665 ;
        RECT 152.560 72.505 152.910 74.665 ;
        RECT 153.390 72.505 153.740 74.665 ;
        RECT 154.220 72.505 154.570 74.665 ;
        RECT 155.050 72.505 155.400 74.665 ;
        RECT 155.880 72.505 156.230 74.665 ;
        RECT 156.710 72.505 157.060 74.665 ;
        RECT 157.540 72.505 157.890 74.665 ;
        RECT 158.370 72.505 158.720 74.665 ;
        RECT 159.200 72.505 159.550 74.665 ;
        RECT 160.030 72.505 160.380 74.665 ;
        RECT 160.860 72.505 161.210 74.665 ;
        RECT 161.690 72.505 162.040 74.665 ;
        RECT 162.520 72.505 162.870 74.665 ;
        RECT 163.350 72.505 163.700 74.665 ;
        RECT 164.180 72.505 164.530 74.665 ;
        RECT 165.010 72.505 165.360 74.665 ;
        RECT 165.840 72.505 166.190 74.665 ;
        RECT 166.670 72.505 167.020 74.665 ;
        RECT 167.500 72.505 167.850 74.665 ;
        RECT 168.330 72.505 168.680 74.665 ;
        RECT 169.160 72.505 169.510 74.665 ;
        RECT 169.990 72.505 170.340 74.665 ;
        RECT 170.820 72.505 171.170 74.665 ;
        RECT 171.650 72.505 172.000 74.665 ;
        RECT 172.480 72.505 172.830 74.665 ;
        RECT 173.310 72.505 173.660 74.665 ;
        RECT 174.140 72.505 174.490 74.665 ;
        RECT 174.970 72.505 175.320 74.665 ;
        RECT 175.800 72.505 176.150 74.665 ;
        RECT 176.630 72.505 176.980 74.665 ;
        RECT 177.460 72.505 177.810 74.665 ;
        RECT 178.290 72.505 178.640 74.665 ;
        RECT 179.120 72.505 179.470 74.665 ;
        RECT 179.950 72.505 180.300 74.665 ;
        RECT 180.780 72.505 181.130 74.665 ;
        RECT 181.610 72.505 181.960 74.665 ;
        RECT 182.440 72.505 182.790 74.665 ;
        RECT 183.270 72.505 183.620 74.665 ;
        RECT 184.100 72.505 184.450 74.665 ;
        RECT 184.930 72.505 185.280 74.665 ;
        RECT 185.760 72.505 186.110 74.665 ;
        RECT 186.590 72.505 186.940 74.665 ;
        RECT 187.420 72.505 187.770 74.665 ;
        RECT 188.250 72.505 188.600 74.665 ;
        RECT 189.080 72.505 189.430 74.665 ;
        RECT 189.910 72.505 190.260 74.665 ;
        RECT 190.740 72.505 191.090 74.665 ;
        RECT 191.570 72.505 191.920 74.665 ;
        RECT 192.400 72.505 192.750 74.665 ;
        RECT 193.230 72.505 193.580 74.665 ;
        RECT 194.060 72.505 194.410 74.665 ;
        RECT 194.890 72.505 195.240 74.665 ;
        RECT 195.720 72.505 196.070 74.665 ;
        RECT 196.550 72.505 196.900 74.665 ;
        RECT 197.380 72.505 197.730 74.665 ;
        RECT 198.210 72.505 198.560 74.665 ;
        RECT 199.040 72.505 199.390 74.665 ;
        RECT 199.870 72.505 200.220 74.665 ;
        RECT 200.700 72.505 201.050 74.665 ;
        RECT 201.530 72.505 201.880 74.665 ;
        RECT 202.360 72.505 202.710 74.665 ;
        RECT 203.190 72.505 203.540 74.665 ;
        RECT 204.020 72.505 204.370 74.665 ;
        RECT 204.850 72.505 205.200 74.665 ;
        RECT 205.680 72.505 206.030 74.665 ;
        RECT 206.510 72.505 206.860 74.665 ;
        RECT 207.340 72.505 207.690 74.665 ;
        RECT 208.170 72.505 208.520 74.665 ;
        RECT 209.000 72.505 209.350 74.665 ;
        RECT 209.830 72.505 210.180 74.665 ;
        RECT 210.660 72.505 211.010 74.665 ;
        RECT 211.490 72.505 211.840 74.665 ;
        RECT 212.320 71.900 212.675 75.145 ;
        RECT 215.625 71.900 228.050 75.945 ;
        RECT 97.780 68.505 98.130 70.665 ;
        RECT 98.610 68.505 98.960 70.665 ;
        RECT 99.440 68.505 99.790 70.665 ;
        RECT 100.270 68.505 100.620 70.665 ;
        RECT 101.100 68.505 101.450 70.665 ;
        RECT 101.930 68.505 102.280 70.665 ;
        RECT 102.760 68.505 103.110 70.665 ;
        RECT 103.590 68.505 103.940 70.665 ;
        RECT 104.420 68.505 104.770 70.665 ;
        RECT 105.250 68.505 105.600 70.665 ;
        RECT 106.080 68.505 106.430 70.665 ;
        RECT 106.910 68.505 107.260 70.665 ;
        RECT 107.740 68.505 108.090 70.665 ;
        RECT 108.570 68.505 108.920 70.665 ;
        RECT 109.400 68.505 109.750 70.665 ;
        RECT 110.230 68.505 110.580 70.665 ;
        RECT 111.060 68.505 111.410 70.665 ;
        RECT 111.890 68.505 112.240 70.665 ;
        RECT 112.720 68.505 113.070 70.665 ;
        RECT 113.550 68.505 113.900 70.665 ;
        RECT 114.380 68.505 114.730 70.665 ;
        RECT 115.210 68.505 115.560 70.665 ;
        RECT 116.040 68.505 116.390 70.665 ;
        RECT 116.870 68.505 117.220 70.665 ;
        RECT 117.700 68.505 118.050 70.665 ;
        RECT 118.530 68.505 118.880 70.665 ;
        RECT 119.360 68.505 119.710 70.665 ;
        RECT 120.190 68.505 120.540 70.665 ;
        RECT 121.020 68.505 121.370 70.665 ;
        RECT 121.850 68.505 122.200 70.665 ;
        RECT 122.680 68.505 123.030 70.665 ;
        RECT 123.510 68.505 123.860 70.665 ;
        RECT 124.340 68.505 124.690 70.665 ;
        RECT 125.170 68.505 125.520 70.665 ;
        RECT 126.000 68.505 126.350 70.665 ;
        RECT 126.830 68.505 127.180 70.665 ;
        RECT 127.660 68.505 128.010 70.665 ;
        RECT 128.490 68.505 128.840 70.665 ;
        RECT 129.320 68.505 129.670 70.665 ;
        RECT 130.150 68.505 130.500 70.665 ;
        RECT 130.980 68.505 131.330 70.665 ;
        RECT 131.810 68.505 132.160 70.665 ;
        RECT 132.640 68.505 132.990 70.665 ;
        RECT 133.470 68.505 133.820 70.665 ;
        RECT 134.300 68.505 134.650 70.665 ;
        RECT 135.130 68.505 135.480 70.665 ;
        RECT 135.960 68.505 136.310 70.665 ;
        RECT 136.790 68.505 137.140 70.665 ;
        RECT 137.620 68.505 137.970 70.665 ;
        RECT 138.450 68.505 138.800 70.665 ;
        RECT 139.280 68.505 139.630 70.665 ;
        RECT 140.110 68.505 140.460 70.665 ;
        RECT 140.940 68.505 141.290 70.665 ;
        RECT 141.770 68.505 142.120 70.665 ;
        RECT 142.600 68.505 142.950 70.665 ;
        RECT 143.430 68.505 143.780 70.665 ;
        RECT 144.260 68.505 144.610 70.665 ;
        RECT 145.090 68.505 145.440 70.665 ;
        RECT 145.920 68.505 146.270 70.665 ;
        RECT 146.750 68.505 147.100 70.665 ;
        RECT 147.580 68.505 147.930 70.665 ;
        RECT 148.410 68.505 148.760 70.665 ;
        RECT 149.240 68.505 149.590 70.665 ;
        RECT 150.070 68.505 150.420 70.665 ;
        RECT 150.900 68.505 151.250 70.665 ;
        RECT 151.730 68.505 152.080 70.665 ;
        RECT 152.560 68.505 152.910 70.665 ;
        RECT 153.390 68.505 153.740 70.665 ;
        RECT 154.220 68.505 154.570 70.665 ;
        RECT 155.050 68.505 155.400 70.665 ;
        RECT 155.880 68.505 156.230 70.665 ;
        RECT 156.710 68.505 157.060 70.665 ;
        RECT 157.540 68.505 157.890 70.665 ;
        RECT 158.370 68.505 158.720 70.665 ;
        RECT 159.200 68.505 159.550 70.665 ;
        RECT 160.030 68.505 160.380 70.665 ;
        RECT 160.860 68.505 161.210 70.665 ;
        RECT 161.690 68.505 162.040 70.665 ;
        RECT 162.520 68.505 162.870 70.665 ;
        RECT 163.350 68.505 163.700 70.665 ;
        RECT 164.180 68.505 164.530 70.665 ;
        RECT 165.010 68.505 165.360 70.665 ;
        RECT 165.840 68.505 166.190 70.665 ;
        RECT 166.670 68.505 167.020 70.665 ;
        RECT 167.500 68.505 167.850 70.665 ;
        RECT 168.330 68.505 168.680 70.665 ;
        RECT 169.160 68.505 169.510 70.665 ;
        RECT 169.990 68.505 170.340 70.665 ;
        RECT 170.820 68.505 171.170 70.665 ;
        RECT 171.650 68.505 172.000 70.665 ;
        RECT 172.480 68.505 172.830 70.665 ;
        RECT 173.310 68.505 173.660 70.665 ;
        RECT 174.140 68.505 174.490 70.665 ;
        RECT 174.970 68.505 175.320 70.665 ;
        RECT 175.800 68.505 176.150 70.665 ;
        RECT 176.630 68.505 176.980 70.665 ;
        RECT 177.460 68.505 177.810 70.665 ;
        RECT 178.290 68.505 178.640 70.665 ;
        RECT 179.120 68.505 179.470 70.665 ;
        RECT 179.950 68.505 180.300 70.665 ;
        RECT 180.780 68.505 181.130 70.665 ;
        RECT 181.610 68.505 181.960 70.665 ;
        RECT 182.440 68.505 182.790 70.665 ;
        RECT 183.270 68.505 183.620 70.665 ;
        RECT 184.100 68.505 184.450 70.665 ;
        RECT 184.930 68.505 185.280 70.665 ;
        RECT 185.760 68.505 186.110 70.665 ;
        RECT 186.590 68.505 186.940 70.665 ;
        RECT 187.420 68.505 187.770 70.665 ;
        RECT 188.250 68.505 188.600 70.665 ;
        RECT 189.080 68.505 189.430 70.665 ;
        RECT 189.910 68.505 190.260 70.665 ;
        RECT 190.740 68.505 191.090 70.665 ;
        RECT 191.570 68.505 191.920 70.665 ;
        RECT 192.400 68.505 192.750 70.665 ;
        RECT 193.230 68.505 193.580 70.665 ;
        RECT 194.060 68.505 194.410 70.665 ;
        RECT 194.890 68.505 195.240 70.665 ;
        RECT 195.720 68.505 196.070 70.665 ;
        RECT 196.550 68.505 196.900 70.665 ;
        RECT 197.380 68.505 197.730 70.665 ;
        RECT 198.210 68.505 198.560 70.665 ;
        RECT 199.040 68.505 199.390 70.665 ;
        RECT 199.870 68.505 200.220 70.665 ;
        RECT 200.700 68.505 201.050 70.665 ;
        RECT 201.530 68.505 201.880 70.665 ;
        RECT 202.360 68.505 202.710 70.665 ;
        RECT 203.190 68.505 203.540 70.665 ;
        RECT 204.020 68.505 204.370 70.665 ;
        RECT 204.850 68.505 205.200 70.665 ;
        RECT 205.680 68.505 206.030 70.665 ;
        RECT 206.510 68.505 206.860 70.665 ;
        RECT 207.340 68.505 207.690 70.665 ;
        RECT 208.170 68.505 208.520 70.665 ;
        RECT 209.000 68.505 209.350 70.665 ;
        RECT 209.830 68.505 210.180 70.665 ;
        RECT 210.660 68.505 211.010 70.665 ;
        RECT 211.490 68.505 211.840 70.665 ;
        RECT 212.320 69.900 228.050 71.900 ;
        RECT 231.050 75.350 233.700 75.355 ;
        RECT 231.050 75.000 254.955 75.350 ;
        RECT 231.050 70.510 231.425 75.000 ;
        RECT 233.325 74.995 254.955 75.000 ;
        RECT 233.325 74.990 249.805 74.995 ;
        RECT 231.950 74.455 232.800 74.830 ;
        RECT 231.810 71.235 231.980 74.275 ;
        RECT 232.290 71.235 232.460 74.275 ;
        RECT 232.770 71.235 232.940 74.275 ;
        RECT 233.325 74.250 236.000 74.990 ;
        RECT 236.270 74.470 236.795 74.795 ;
        RECT 238.095 74.470 238.620 74.795 ;
        RECT 236.400 74.250 236.570 74.265 ;
        RECT 236.880 74.250 237.050 74.265 ;
        RECT 233.325 71.225 237.075 74.250 ;
        RECT 237.360 71.225 237.530 74.265 ;
        RECT 237.840 74.250 238.010 74.265 ;
        RECT 238.320 74.250 238.490 74.265 ;
        RECT 238.890 74.250 240.600 74.990 ;
        RECT 242.570 74.470 242.945 74.795 ;
        RECT 241.000 74.250 241.170 74.265 ;
        RECT 241.480 74.250 241.650 74.265 ;
        RECT 237.825 71.225 241.675 74.250 ;
        RECT 241.960 71.225 242.130 74.265 ;
        RECT 242.440 74.250 242.610 74.265 ;
        RECT 242.920 74.250 243.090 74.265 ;
        RECT 243.490 74.250 245.200 74.990 ;
        RECT 245.470 74.470 245.995 74.795 ;
        RECT 247.295 74.470 247.820 74.795 ;
        RECT 248.090 74.275 249.805 74.990 ;
        RECT 250.080 74.475 250.580 74.800 ;
        RECT 253.830 74.475 254.330 74.800 ;
        RECT 254.605 74.275 254.955 74.995 ;
        RECT 245.600 74.250 245.770 74.265 ;
        RECT 246.080 74.250 246.250 74.265 ;
        RECT 242.425 71.225 246.275 74.250 ;
        RECT 246.560 71.225 246.730 74.265 ;
        RECT 247.040 74.250 247.210 74.265 ;
        RECT 247.520 74.250 247.690 74.265 ;
        RECT 248.090 74.250 250.875 74.275 ;
        RECT 247.025 71.225 250.875 74.250 ;
        RECT 251.160 71.230 251.330 74.270 ;
        RECT 251.640 71.230 251.810 74.270 ;
        RECT 252.120 71.230 252.290 74.270 ;
        RECT 252.600 71.230 252.770 74.270 ;
        RECT 253.080 71.230 253.250 74.270 ;
        RECT 253.525 71.225 254.955 74.275 ;
        RECT 256.625 74.100 256.975 78.590 ;
        RECT 257.540 78.045 259.290 78.420 ;
        RECT 268.590 78.045 270.340 78.420 ;
        RECT 257.375 74.825 257.545 77.865 ;
        RECT 257.855 74.825 258.025 77.865 ;
        RECT 258.335 74.825 258.505 77.865 ;
        RECT 258.815 74.825 258.985 77.865 ;
        RECT 259.295 74.825 259.465 77.865 ;
        RECT 259.775 74.825 259.945 77.865 ;
        RECT 260.255 74.825 260.425 77.865 ;
        RECT 260.735 74.825 260.905 77.865 ;
        RECT 261.215 74.825 261.385 77.865 ;
        RECT 261.695 74.825 261.865 77.865 ;
        RECT 262.175 74.825 262.345 77.865 ;
        RECT 262.655 74.825 262.825 77.865 ;
        RECT 263.135 74.825 263.305 77.865 ;
        RECT 263.615 74.825 263.785 77.865 ;
        RECT 264.095 74.825 264.265 77.865 ;
        RECT 264.575 74.825 264.745 77.865 ;
        RECT 265.055 74.825 265.225 77.865 ;
        RECT 265.535 74.825 265.705 77.865 ;
        RECT 266.015 74.825 266.185 77.865 ;
        RECT 266.495 74.825 266.665 77.865 ;
        RECT 266.975 74.825 267.145 77.865 ;
        RECT 267.455 74.825 267.625 77.865 ;
        RECT 267.935 74.825 268.105 77.865 ;
        RECT 268.415 74.825 268.585 77.865 ;
        RECT 268.895 74.825 269.065 77.865 ;
        RECT 269.375 74.825 269.545 77.865 ;
        RECT 269.855 74.825 270.025 77.865 ;
        RECT 270.335 74.825 270.505 77.865 ;
        RECT 259.465 74.270 268.415 74.645 ;
        RECT 270.900 74.100 271.250 78.590 ;
        RECT 256.625 73.750 271.250 74.100 ;
        RECT 233.325 70.510 236.000 71.225 ;
        RECT 237.045 70.670 237.845 71.045 ;
        RECT 231.050 70.500 236.000 70.510 ;
        RECT 238.890 70.500 240.600 71.225 ;
        RECT 242.095 70.670 242.470 71.045 ;
        RECT 243.490 70.500 245.200 71.225 ;
        RECT 246.245 70.670 247.045 71.045 ;
        RECT 248.090 70.505 249.805 71.225 ;
        RECT 250.830 70.675 253.580 71.050 ;
        RECT 254.605 70.505 254.955 71.225 ;
        RECT 248.090 70.500 254.955 70.505 ;
        RECT 231.050 70.155 254.955 70.500 ;
        RECT 233.325 70.150 254.955 70.155 ;
        RECT 256.625 73.150 271.250 73.500 ;
        RECT 256.625 70.750 256.975 73.150 ;
        RECT 257.540 72.650 259.290 72.975 ;
        RECT 268.590 72.650 270.340 72.975 ;
        RECT 257.375 71.430 257.545 72.470 ;
        RECT 257.855 71.430 258.025 72.470 ;
        RECT 258.335 71.430 258.505 72.470 ;
        RECT 258.815 71.430 258.985 72.470 ;
        RECT 259.295 71.430 259.465 72.470 ;
        RECT 259.775 71.430 259.945 72.470 ;
        RECT 260.255 71.430 260.425 72.470 ;
        RECT 260.735 71.430 260.905 72.470 ;
        RECT 261.215 71.430 261.385 72.470 ;
        RECT 261.695 71.430 261.865 72.470 ;
        RECT 262.175 71.430 262.345 72.470 ;
        RECT 262.655 71.430 262.825 72.470 ;
        RECT 263.135 71.430 263.305 72.470 ;
        RECT 263.615 71.430 263.785 72.470 ;
        RECT 264.095 71.430 264.265 72.470 ;
        RECT 264.575 71.430 264.745 72.470 ;
        RECT 265.055 71.430 265.225 72.470 ;
        RECT 265.535 71.430 265.705 72.470 ;
        RECT 266.015 71.430 266.185 72.470 ;
        RECT 266.495 71.430 266.665 72.470 ;
        RECT 266.975 71.430 267.145 72.470 ;
        RECT 267.455 71.430 267.625 72.470 ;
        RECT 267.935 71.430 268.105 72.470 ;
        RECT 268.415 71.430 268.585 72.470 ;
        RECT 268.895 71.430 269.065 72.470 ;
        RECT 269.375 71.430 269.545 72.470 ;
        RECT 269.855 71.430 270.025 72.470 ;
        RECT 270.335 71.430 270.505 72.470 ;
        RECT 259.465 70.925 268.415 71.250 ;
        RECT 270.900 70.750 271.250 73.150 ;
        RECT 235.645 70.145 239.245 70.150 ;
        RECT 240.245 70.145 243.845 70.150 ;
        RECT 244.845 70.145 248.445 70.150 ;
        RECT 212.320 69.875 254.955 69.900 ;
        RECT 256.625 69.875 271.250 70.750 ;
        RECT 212.320 69.550 271.250 69.875 ;
        RECT 212.320 68.025 231.425 69.550 ;
        RECT 233.325 68.875 236.005 69.550 ;
        RECT 237.050 69.050 237.850 69.375 ;
        RECT 238.895 68.875 240.605 69.550 ;
        RECT 242.100 69.050 242.475 69.375 ;
        RECT 243.495 68.875 245.205 69.550 ;
        RECT 246.250 69.050 247.050 69.375 ;
        RECT 248.095 68.875 249.805 69.550 ;
        RECT 250.830 69.050 253.580 69.375 ;
        RECT 254.605 68.875 271.250 69.550 ;
        RECT 75.275 67.150 231.425 68.025 ;
        RECT 231.810 67.830 231.980 68.870 ;
        RECT 232.290 67.830 232.460 68.870 ;
        RECT 232.770 67.830 232.940 68.870 ;
        RECT 233.325 67.825 237.075 68.875 ;
        RECT 237.365 67.830 237.535 68.870 ;
        RECT 237.825 67.825 241.675 68.875 ;
        RECT 241.965 67.830 242.135 68.870 ;
        RECT 242.425 67.825 246.275 68.875 ;
        RECT 246.565 67.830 246.735 68.870 ;
        RECT 247.025 67.825 250.875 68.875 ;
        RECT 251.160 67.830 251.330 68.870 ;
        RECT 251.640 67.830 251.810 68.870 ;
        RECT 252.120 67.830 252.290 68.870 ;
        RECT 252.600 67.830 252.770 68.870 ;
        RECT 253.080 67.830 253.250 68.870 ;
        RECT 253.525 67.825 271.250 68.875 ;
        RECT 231.950 67.325 232.800 67.650 ;
        RECT 233.325 67.150 236.005 67.825 ;
        RECT 236.275 67.325 236.800 67.650 ;
        RECT 238.100 67.325 238.625 67.650 ;
        RECT 238.895 67.150 240.605 67.825 ;
        RECT 242.575 67.325 242.950 67.650 ;
        RECT 243.495 67.150 245.205 67.825 ;
        RECT 245.475 67.325 246.000 67.650 ;
        RECT 247.300 67.325 247.825 67.650 ;
        RECT 248.095 67.150 249.805 67.825 ;
        RECT 250.080 67.325 250.580 67.650 ;
        RECT 253.830 67.325 254.330 67.650 ;
        RECT 254.605 67.150 271.250 67.825 ;
        RECT 75.275 65.950 271.250 67.150 ;
      LAYER met1 ;
        RECT 138.275 213.850 237.100 214.450 ;
        RECT 135.525 210.575 233.850 211.175 ;
        RECT 132.775 207.300 230.600 207.900 ;
        RECT 130.000 204.050 227.350 204.650 ;
        RECT 226.750 161.675 227.350 204.050 ;
        RECT 226.750 161.075 229.275 161.675 ;
        RECT 75.275 157.875 228.050 159.850 ;
        RECT 75.275 154.000 97.300 157.875 ;
        RECT 97.830 157.325 98.080 157.360 ;
        RECT 98.660 157.325 98.910 157.360 ;
        RECT 99.490 157.325 99.740 157.360 ;
        RECT 100.320 157.325 100.570 157.360 ;
        RECT 101.150 157.325 101.400 157.360 ;
        RECT 101.980 157.325 102.230 157.360 ;
        RECT 102.810 157.325 103.060 157.360 ;
        RECT 103.640 157.325 103.890 157.360 ;
        RECT 104.470 157.325 104.720 157.360 ;
        RECT 105.300 157.325 105.550 157.360 ;
        RECT 106.130 157.325 106.380 157.360 ;
        RECT 106.960 157.325 107.210 157.360 ;
        RECT 107.790 157.325 108.040 157.360 ;
        RECT 108.620 157.325 108.870 157.360 ;
        RECT 109.450 157.325 109.700 157.360 ;
        RECT 110.280 157.325 110.530 157.360 ;
        RECT 111.110 157.325 111.360 157.360 ;
        RECT 111.940 157.325 112.190 157.360 ;
        RECT 112.770 157.325 113.020 157.360 ;
        RECT 113.600 157.325 113.850 157.360 ;
        RECT 114.430 157.325 114.680 157.360 ;
        RECT 115.260 157.325 115.510 157.360 ;
        RECT 116.090 157.325 116.340 157.360 ;
        RECT 116.920 157.325 117.170 157.360 ;
        RECT 117.750 157.325 118.000 157.360 ;
        RECT 118.580 157.325 118.830 157.360 ;
        RECT 119.410 157.325 119.660 157.360 ;
        RECT 120.240 157.325 120.490 157.360 ;
        RECT 121.070 157.325 121.320 157.360 ;
        RECT 121.900 157.325 122.150 157.360 ;
        RECT 122.730 157.325 122.980 157.360 ;
        RECT 123.560 157.325 123.810 157.360 ;
        RECT 124.390 157.325 124.640 157.360 ;
        RECT 125.220 157.325 125.470 157.360 ;
        RECT 126.050 157.325 126.300 157.360 ;
        RECT 126.880 157.325 127.130 157.360 ;
        RECT 97.825 155.300 98.925 157.325 ;
        RECT 99.475 155.300 100.575 157.325 ;
        RECT 101.150 155.300 102.250 157.325 ;
        RECT 102.800 155.300 103.900 157.325 ;
        RECT 104.470 155.300 105.575 157.325 ;
        RECT 106.125 155.300 107.225 157.325 ;
        RECT 107.790 155.300 108.900 157.325 ;
        RECT 109.450 155.300 110.550 157.325 ;
        RECT 111.100 155.300 112.200 157.325 ;
        RECT 112.770 155.300 113.875 157.325 ;
        RECT 114.425 155.300 115.525 157.325 ;
        RECT 116.090 155.300 117.200 157.325 ;
        RECT 117.750 155.300 118.850 157.325 ;
        RECT 119.400 155.300 120.500 157.325 ;
        RECT 121.070 155.300 122.175 157.325 ;
        RECT 122.725 155.300 123.825 157.325 ;
        RECT 124.390 155.300 125.500 157.325 ;
        RECT 126.050 155.300 127.150 157.325 ;
        RECT 97.830 155.255 98.080 155.300 ;
        RECT 98.660 155.255 98.910 155.300 ;
        RECT 99.490 155.255 99.740 155.300 ;
        RECT 100.320 155.255 100.570 155.300 ;
        RECT 101.150 155.255 101.400 155.300 ;
        RECT 101.980 155.255 102.230 155.300 ;
        RECT 102.810 155.255 103.060 155.300 ;
        RECT 103.640 155.255 103.890 155.300 ;
        RECT 104.470 155.255 104.720 155.300 ;
        RECT 105.300 155.255 105.550 155.300 ;
        RECT 106.130 155.255 106.380 155.300 ;
        RECT 106.960 155.255 107.210 155.300 ;
        RECT 107.790 155.255 108.040 155.300 ;
        RECT 108.620 155.255 108.870 155.300 ;
        RECT 109.450 155.255 109.700 155.300 ;
        RECT 110.280 155.255 110.530 155.300 ;
        RECT 111.110 155.255 111.360 155.300 ;
        RECT 111.940 155.255 112.190 155.300 ;
        RECT 112.770 155.255 113.020 155.300 ;
        RECT 113.600 155.255 113.850 155.300 ;
        RECT 114.430 155.255 114.680 155.300 ;
        RECT 115.260 155.255 115.510 155.300 ;
        RECT 116.090 155.255 116.340 155.300 ;
        RECT 116.920 155.255 117.170 155.300 ;
        RECT 117.750 155.255 118.000 155.300 ;
        RECT 118.580 155.255 118.830 155.300 ;
        RECT 119.410 155.255 119.660 155.300 ;
        RECT 120.240 155.255 120.490 155.300 ;
        RECT 121.070 155.255 121.320 155.300 ;
        RECT 121.900 155.255 122.150 155.300 ;
        RECT 122.730 155.255 122.980 155.300 ;
        RECT 123.560 155.255 123.810 155.300 ;
        RECT 124.390 155.255 124.640 155.300 ;
        RECT 125.220 155.255 125.470 155.300 ;
        RECT 126.050 155.255 126.300 155.300 ;
        RECT 126.880 155.255 127.130 155.300 ;
        RECT 127.675 155.250 128.825 157.375 ;
        RECT 129.370 157.325 129.620 157.360 ;
        RECT 130.200 157.325 130.450 157.360 ;
        RECT 131.030 157.325 131.280 157.360 ;
        RECT 131.860 157.325 132.110 157.360 ;
        RECT 132.690 157.325 132.940 157.360 ;
        RECT 133.520 157.325 133.770 157.360 ;
        RECT 134.350 157.325 134.600 157.360 ;
        RECT 135.180 157.325 135.430 157.360 ;
        RECT 136.010 157.325 136.260 157.360 ;
        RECT 136.840 157.325 137.090 157.360 ;
        RECT 137.670 157.325 137.920 157.360 ;
        RECT 138.500 157.325 138.750 157.360 ;
        RECT 139.330 157.325 139.580 157.360 ;
        RECT 140.160 157.325 140.410 157.360 ;
        RECT 140.990 157.325 141.240 157.360 ;
        RECT 141.820 157.325 142.070 157.360 ;
        RECT 142.650 157.325 142.900 157.360 ;
        RECT 143.480 157.325 143.730 157.360 ;
        RECT 144.310 157.325 144.560 157.360 ;
        RECT 145.140 157.325 145.390 157.360 ;
        RECT 145.970 157.325 146.220 157.360 ;
        RECT 146.800 157.325 147.050 157.360 ;
        RECT 147.630 157.325 147.880 157.360 ;
        RECT 148.460 157.325 148.710 157.360 ;
        RECT 149.290 157.325 149.540 157.360 ;
        RECT 150.120 157.325 150.370 157.360 ;
        RECT 150.950 157.325 151.200 157.360 ;
        RECT 151.780 157.325 152.030 157.360 ;
        RECT 152.610 157.325 152.860 157.360 ;
        RECT 153.440 157.325 153.690 157.360 ;
        RECT 154.270 157.325 154.520 157.360 ;
        RECT 155.100 157.325 155.350 157.360 ;
        RECT 155.930 157.325 156.180 157.360 ;
        RECT 156.760 157.325 157.010 157.360 ;
        RECT 157.590 157.325 157.840 157.360 ;
        RECT 158.420 157.325 158.670 157.360 ;
        RECT 159.250 157.325 159.500 157.360 ;
        RECT 160.080 157.325 160.330 157.360 ;
        RECT 160.910 157.325 161.160 157.360 ;
        RECT 161.740 157.325 161.990 157.360 ;
        RECT 162.570 157.325 162.820 157.360 ;
        RECT 163.400 157.325 163.650 157.360 ;
        RECT 164.230 157.325 164.480 157.360 ;
        RECT 165.060 157.325 165.310 157.360 ;
        RECT 165.890 157.325 166.140 157.360 ;
        RECT 166.720 157.325 166.970 157.360 ;
        RECT 167.550 157.325 167.800 157.360 ;
        RECT 168.380 157.325 168.630 157.360 ;
        RECT 169.210 157.325 169.460 157.360 ;
        RECT 170.040 157.325 170.290 157.360 ;
        RECT 170.870 157.325 171.120 157.360 ;
        RECT 171.700 157.325 171.950 157.360 ;
        RECT 172.530 157.325 172.780 157.360 ;
        RECT 173.360 157.325 173.610 157.360 ;
        RECT 174.190 157.325 174.440 157.360 ;
        RECT 175.020 157.325 175.270 157.360 ;
        RECT 175.850 157.325 176.100 157.360 ;
        RECT 176.680 157.325 176.930 157.360 ;
        RECT 177.510 157.325 177.760 157.360 ;
        RECT 178.340 157.325 178.590 157.360 ;
        RECT 179.170 157.325 179.420 157.360 ;
        RECT 180.000 157.325 180.250 157.360 ;
        RECT 180.830 157.325 181.080 157.360 ;
        RECT 181.660 157.325 181.910 157.360 ;
        RECT 182.490 157.325 182.740 157.360 ;
        RECT 183.320 157.325 183.570 157.360 ;
        RECT 184.150 157.325 184.400 157.360 ;
        RECT 184.980 157.325 185.230 157.360 ;
        RECT 185.810 157.325 186.060 157.360 ;
        RECT 186.640 157.325 186.890 157.360 ;
        RECT 187.470 157.325 187.720 157.360 ;
        RECT 188.300 157.325 188.550 157.360 ;
        RECT 189.130 157.325 189.380 157.360 ;
        RECT 189.960 157.325 190.210 157.360 ;
        RECT 190.790 157.325 191.040 157.360 ;
        RECT 191.620 157.325 191.870 157.360 ;
        RECT 192.450 157.325 192.700 157.360 ;
        RECT 193.280 157.325 193.530 157.360 ;
        RECT 194.110 157.325 194.360 157.360 ;
        RECT 194.940 157.325 195.190 157.360 ;
        RECT 195.770 157.325 196.020 157.360 ;
        RECT 196.600 157.325 196.850 157.360 ;
        RECT 197.430 157.325 197.680 157.360 ;
        RECT 198.260 157.325 198.510 157.360 ;
        RECT 199.090 157.325 199.340 157.360 ;
        RECT 199.920 157.325 200.170 157.360 ;
        RECT 200.750 157.325 201.000 157.360 ;
        RECT 201.580 157.325 201.830 157.360 ;
        RECT 202.410 157.325 202.660 157.360 ;
        RECT 203.240 157.325 203.490 157.360 ;
        RECT 204.070 157.325 204.320 157.360 ;
        RECT 204.900 157.325 205.150 157.360 ;
        RECT 205.730 157.325 205.980 157.360 ;
        RECT 206.560 157.325 206.810 157.360 ;
        RECT 207.390 157.325 207.640 157.360 ;
        RECT 208.220 157.325 208.470 157.360 ;
        RECT 209.050 157.325 209.300 157.360 ;
        RECT 209.880 157.325 210.130 157.360 ;
        RECT 210.710 157.325 210.960 157.360 ;
        RECT 211.540 157.325 211.790 157.360 ;
        RECT 129.370 155.300 130.475 157.325 ;
        RECT 131.025 155.300 132.125 157.325 ;
        RECT 132.690 155.300 133.800 157.325 ;
        RECT 134.350 155.300 135.450 157.325 ;
        RECT 136.000 155.300 137.100 157.325 ;
        RECT 137.670 155.300 138.775 157.325 ;
        RECT 139.325 155.300 140.425 157.325 ;
        RECT 140.990 155.300 142.100 157.325 ;
        RECT 142.650 155.300 143.750 157.325 ;
        RECT 144.300 155.300 145.400 157.325 ;
        RECT 145.950 155.300 147.050 157.325 ;
        RECT 147.625 155.300 148.725 157.325 ;
        RECT 149.290 155.300 150.400 157.325 ;
        RECT 150.950 155.300 152.050 157.325 ;
        RECT 152.600 155.300 153.700 157.325 ;
        RECT 154.270 155.300 155.375 157.325 ;
        RECT 155.925 155.300 157.025 157.325 ;
        RECT 157.575 155.300 158.675 157.325 ;
        RECT 159.250 155.300 160.350 157.325 ;
        RECT 160.900 155.300 162.000 157.325 ;
        RECT 162.570 155.300 163.675 157.325 ;
        RECT 164.225 155.300 165.325 157.325 ;
        RECT 165.890 155.300 167.000 157.325 ;
        RECT 167.550 155.300 168.650 157.325 ;
        RECT 169.200 155.300 170.300 157.325 ;
        RECT 170.870 155.300 171.975 157.325 ;
        RECT 172.525 155.300 173.625 157.325 ;
        RECT 174.190 155.300 175.300 157.325 ;
        RECT 175.850 155.300 176.950 157.325 ;
        RECT 177.500 155.300 178.600 157.325 ;
        RECT 179.170 155.300 180.275 157.325 ;
        RECT 180.825 155.300 181.925 157.325 ;
        RECT 182.490 155.300 183.600 157.325 ;
        RECT 184.150 155.300 185.250 157.325 ;
        RECT 185.800 155.300 186.900 157.325 ;
        RECT 187.470 155.300 188.575 157.325 ;
        RECT 189.125 155.300 190.225 157.325 ;
        RECT 190.790 155.300 191.900 157.325 ;
        RECT 192.450 155.300 193.550 157.325 ;
        RECT 194.100 155.300 195.200 157.325 ;
        RECT 195.770 155.300 196.875 157.325 ;
        RECT 197.425 155.300 198.525 157.325 ;
        RECT 199.090 155.300 200.200 157.325 ;
        RECT 200.750 155.300 201.850 157.325 ;
        RECT 202.400 155.300 203.500 157.325 ;
        RECT 204.070 155.300 205.175 157.325 ;
        RECT 205.725 155.300 206.825 157.325 ;
        RECT 207.390 155.300 208.500 157.325 ;
        RECT 209.050 155.300 210.150 157.325 ;
        RECT 210.700 155.300 211.800 157.325 ;
        RECT 129.370 155.255 129.620 155.300 ;
        RECT 130.200 155.255 130.450 155.300 ;
        RECT 131.030 155.255 131.280 155.300 ;
        RECT 131.860 155.255 132.110 155.300 ;
        RECT 132.690 155.255 132.940 155.300 ;
        RECT 133.520 155.255 133.770 155.300 ;
        RECT 134.350 155.255 134.600 155.300 ;
        RECT 135.180 155.255 135.430 155.300 ;
        RECT 136.010 155.255 136.260 155.300 ;
        RECT 136.840 155.255 137.090 155.300 ;
        RECT 137.670 155.255 137.920 155.300 ;
        RECT 138.500 155.255 138.750 155.300 ;
        RECT 139.330 155.255 139.580 155.300 ;
        RECT 140.160 155.255 140.410 155.300 ;
        RECT 140.990 155.255 141.240 155.300 ;
        RECT 141.820 155.255 142.070 155.300 ;
        RECT 142.650 155.255 142.900 155.300 ;
        RECT 143.480 155.255 143.730 155.300 ;
        RECT 144.310 155.255 144.560 155.300 ;
        RECT 145.140 155.255 145.390 155.300 ;
        RECT 145.970 155.255 146.220 155.300 ;
        RECT 146.800 155.255 147.050 155.300 ;
        RECT 147.630 155.255 147.880 155.300 ;
        RECT 148.460 155.255 148.710 155.300 ;
        RECT 149.290 155.255 149.540 155.300 ;
        RECT 150.120 155.255 150.370 155.300 ;
        RECT 150.950 155.255 151.200 155.300 ;
        RECT 151.780 155.255 152.030 155.300 ;
        RECT 152.610 155.255 152.860 155.300 ;
        RECT 153.440 155.255 153.690 155.300 ;
        RECT 154.270 155.255 154.520 155.300 ;
        RECT 155.100 155.255 155.350 155.300 ;
        RECT 155.930 155.255 156.180 155.300 ;
        RECT 156.760 155.255 157.010 155.300 ;
        RECT 157.590 155.255 157.840 155.300 ;
        RECT 158.420 155.255 158.670 155.300 ;
        RECT 159.250 155.255 159.500 155.300 ;
        RECT 160.080 155.255 160.330 155.300 ;
        RECT 160.910 155.255 161.160 155.300 ;
        RECT 161.740 155.255 161.990 155.300 ;
        RECT 162.570 155.255 162.820 155.300 ;
        RECT 163.400 155.255 163.650 155.300 ;
        RECT 164.230 155.255 164.480 155.300 ;
        RECT 165.060 155.255 165.310 155.300 ;
        RECT 165.890 155.255 166.140 155.300 ;
        RECT 166.720 155.255 166.970 155.300 ;
        RECT 167.550 155.255 167.800 155.300 ;
        RECT 168.380 155.255 168.630 155.300 ;
        RECT 169.210 155.255 169.460 155.300 ;
        RECT 170.040 155.255 170.290 155.300 ;
        RECT 170.870 155.255 171.120 155.300 ;
        RECT 171.700 155.255 171.950 155.300 ;
        RECT 172.530 155.255 172.780 155.300 ;
        RECT 173.360 155.255 173.610 155.300 ;
        RECT 174.190 155.255 174.440 155.300 ;
        RECT 175.020 155.255 175.270 155.300 ;
        RECT 175.850 155.255 176.100 155.300 ;
        RECT 176.680 155.255 176.930 155.300 ;
        RECT 177.510 155.255 177.760 155.300 ;
        RECT 178.340 155.255 178.590 155.300 ;
        RECT 179.170 155.255 179.420 155.300 ;
        RECT 180.000 155.255 180.250 155.300 ;
        RECT 180.830 155.255 181.080 155.300 ;
        RECT 181.660 155.255 181.910 155.300 ;
        RECT 182.490 155.255 182.740 155.300 ;
        RECT 183.320 155.255 183.570 155.300 ;
        RECT 184.150 155.255 184.400 155.300 ;
        RECT 184.980 155.255 185.230 155.300 ;
        RECT 185.810 155.255 186.060 155.300 ;
        RECT 186.640 155.255 186.890 155.300 ;
        RECT 187.470 155.255 187.720 155.300 ;
        RECT 188.300 155.255 188.550 155.300 ;
        RECT 189.130 155.255 189.380 155.300 ;
        RECT 189.960 155.255 190.210 155.300 ;
        RECT 190.790 155.255 191.040 155.300 ;
        RECT 191.620 155.255 191.870 155.300 ;
        RECT 192.450 155.255 192.700 155.300 ;
        RECT 193.280 155.255 193.530 155.300 ;
        RECT 194.110 155.255 194.360 155.300 ;
        RECT 194.940 155.255 195.190 155.300 ;
        RECT 195.770 155.255 196.020 155.300 ;
        RECT 196.600 155.255 196.850 155.300 ;
        RECT 197.430 155.255 197.680 155.300 ;
        RECT 198.260 155.255 198.510 155.300 ;
        RECT 199.090 155.255 199.340 155.300 ;
        RECT 199.920 155.255 200.170 155.300 ;
        RECT 200.750 155.255 201.000 155.300 ;
        RECT 201.580 155.255 201.830 155.300 ;
        RECT 202.410 155.255 202.660 155.300 ;
        RECT 203.240 155.255 203.490 155.300 ;
        RECT 204.070 155.255 204.320 155.300 ;
        RECT 204.900 155.255 205.150 155.300 ;
        RECT 205.730 155.255 205.980 155.300 ;
        RECT 206.560 155.255 206.810 155.300 ;
        RECT 207.390 155.255 207.640 155.300 ;
        RECT 208.220 155.255 208.470 155.300 ;
        RECT 209.050 155.255 209.300 155.300 ;
        RECT 209.880 155.255 210.130 155.300 ;
        RECT 210.710 155.255 210.960 155.300 ;
        RECT 211.540 155.255 211.790 155.300 ;
        RECT 212.325 154.000 228.050 157.875 ;
        RECT 97.830 153.325 98.080 153.365 ;
        RECT 98.660 153.325 98.910 153.365 ;
        RECT 99.490 153.325 99.740 153.365 ;
        RECT 100.320 153.325 100.570 153.365 ;
        RECT 101.150 153.325 101.400 153.365 ;
        RECT 101.980 153.325 102.230 153.365 ;
        RECT 102.810 153.325 103.060 153.365 ;
        RECT 103.640 153.325 103.890 153.365 ;
        RECT 104.470 153.325 104.720 153.365 ;
        RECT 105.300 153.325 105.550 153.365 ;
        RECT 106.130 153.325 106.380 153.365 ;
        RECT 106.960 153.325 107.210 153.365 ;
        RECT 107.790 153.325 108.040 153.365 ;
        RECT 108.620 153.325 108.870 153.365 ;
        RECT 109.450 153.325 109.700 153.365 ;
        RECT 110.280 153.325 110.530 153.365 ;
        RECT 111.110 153.325 111.360 153.365 ;
        RECT 111.940 153.350 112.190 153.365 ;
        RECT 112.770 153.350 113.020 153.365 ;
        RECT 39.400 151.300 98.100 153.325 ;
        RECT 98.650 151.300 99.750 153.325 ;
        RECT 100.300 151.300 101.425 153.325 ;
        RECT 101.975 151.300 103.075 153.325 ;
        RECT 103.625 151.300 104.725 153.325 ;
        RECT 105.300 151.300 106.400 153.325 ;
        RECT 106.950 151.300 108.050 153.325 ;
        RECT 108.600 151.300 109.700 153.325 ;
        RECT 110.275 151.300 111.375 153.325 ;
        RECT 39.400 7.575 41.425 151.300 ;
        RECT 97.830 151.260 98.080 151.300 ;
        RECT 98.660 151.260 98.910 151.300 ;
        RECT 99.490 151.260 99.740 151.300 ;
        RECT 100.320 151.260 100.570 151.300 ;
        RECT 101.150 151.260 101.400 151.300 ;
        RECT 101.980 151.260 102.230 151.300 ;
        RECT 102.810 151.260 103.060 151.300 ;
        RECT 103.640 151.260 103.890 151.300 ;
        RECT 104.470 151.260 104.720 151.300 ;
        RECT 105.300 151.260 105.550 151.300 ;
        RECT 106.130 151.260 106.380 151.300 ;
        RECT 106.960 151.260 107.210 151.300 ;
        RECT 107.790 151.260 108.040 151.300 ;
        RECT 108.620 151.260 108.870 151.300 ;
        RECT 109.450 151.260 109.700 151.300 ;
        RECT 110.280 151.260 110.530 151.300 ;
        RECT 111.110 151.260 111.360 151.300 ;
        RECT 111.925 151.125 113.050 153.350 ;
        RECT 113.600 153.325 113.850 153.365 ;
        RECT 114.430 153.325 114.680 153.365 ;
        RECT 115.260 153.325 115.510 153.365 ;
        RECT 116.090 153.325 116.340 153.365 ;
        RECT 116.920 153.325 117.170 153.365 ;
        RECT 117.750 153.325 118.000 153.365 ;
        RECT 118.580 153.325 118.830 153.365 ;
        RECT 119.410 153.325 119.660 153.365 ;
        RECT 120.240 153.325 120.490 153.365 ;
        RECT 121.070 153.325 121.320 153.365 ;
        RECT 121.900 153.325 122.150 153.365 ;
        RECT 122.730 153.325 122.980 153.365 ;
        RECT 123.560 153.325 123.810 153.365 ;
        RECT 124.390 153.325 124.640 153.365 ;
        RECT 125.220 153.325 125.470 153.365 ;
        RECT 126.050 153.325 126.300 153.365 ;
        RECT 126.880 153.325 127.130 153.365 ;
        RECT 127.710 153.325 127.960 153.365 ;
        RECT 128.540 153.325 128.790 153.365 ;
        RECT 129.370 153.325 129.620 153.365 ;
        RECT 130.200 153.325 130.450 153.365 ;
        RECT 131.030 153.325 131.280 153.365 ;
        RECT 131.860 153.325 132.110 153.365 ;
        RECT 132.690 153.325 132.940 153.365 ;
        RECT 133.520 153.325 133.770 153.365 ;
        RECT 134.350 153.325 134.600 153.365 ;
        RECT 135.180 153.325 135.430 153.365 ;
        RECT 136.010 153.325 136.260 153.365 ;
        RECT 136.840 153.325 137.090 153.365 ;
        RECT 137.670 153.325 137.920 153.365 ;
        RECT 138.500 153.325 138.750 153.365 ;
        RECT 139.330 153.325 139.580 153.365 ;
        RECT 140.160 153.325 140.410 153.365 ;
        RECT 140.990 153.325 141.240 153.365 ;
        RECT 141.820 153.325 142.070 153.365 ;
        RECT 142.650 153.325 142.900 153.365 ;
        RECT 143.480 153.325 143.730 153.365 ;
        RECT 144.310 153.325 144.560 153.365 ;
        RECT 145.140 153.325 145.390 153.365 ;
        RECT 145.970 153.325 146.220 153.365 ;
        RECT 146.800 153.325 147.050 153.365 ;
        RECT 147.630 153.325 147.880 153.365 ;
        RECT 148.460 153.325 148.710 153.365 ;
        RECT 149.290 153.325 149.540 153.365 ;
        RECT 150.120 153.325 150.370 153.365 ;
        RECT 150.950 153.325 151.200 153.365 ;
        RECT 151.780 153.325 152.030 153.365 ;
        RECT 152.610 153.325 152.860 153.365 ;
        RECT 153.440 153.325 153.690 153.365 ;
        RECT 154.270 153.325 154.520 153.365 ;
        RECT 155.100 153.325 155.350 153.365 ;
        RECT 155.930 153.325 156.180 153.365 ;
        RECT 156.760 153.325 157.010 153.365 ;
        RECT 157.590 153.325 157.840 153.365 ;
        RECT 158.420 153.325 158.670 153.365 ;
        RECT 159.250 153.325 159.500 153.365 ;
        RECT 160.080 153.325 160.330 153.365 ;
        RECT 160.910 153.325 161.160 153.365 ;
        RECT 161.740 153.325 161.990 153.365 ;
        RECT 162.570 153.325 162.820 153.365 ;
        RECT 163.400 153.325 163.650 153.365 ;
        RECT 164.230 153.325 164.480 153.365 ;
        RECT 165.060 153.325 165.310 153.365 ;
        RECT 165.890 153.325 166.140 153.365 ;
        RECT 166.720 153.325 166.970 153.365 ;
        RECT 167.550 153.325 167.800 153.365 ;
        RECT 168.380 153.325 168.630 153.365 ;
        RECT 169.210 153.325 169.460 153.365 ;
        RECT 170.040 153.325 170.290 153.365 ;
        RECT 170.870 153.325 171.120 153.365 ;
        RECT 171.700 153.325 171.950 153.365 ;
        RECT 172.530 153.325 172.780 153.365 ;
        RECT 173.360 153.325 173.610 153.365 ;
        RECT 174.190 153.325 174.440 153.365 ;
        RECT 175.020 153.325 175.270 153.365 ;
        RECT 175.850 153.325 176.100 153.365 ;
        RECT 176.680 153.325 176.930 153.365 ;
        RECT 177.510 153.325 177.760 153.365 ;
        RECT 178.340 153.325 178.590 153.365 ;
        RECT 179.170 153.325 179.420 153.365 ;
        RECT 113.600 151.300 114.700 153.325 ;
        RECT 115.250 151.300 116.350 153.325 ;
        RECT 116.920 151.300 118.025 153.325 ;
        RECT 118.575 151.300 119.675 153.325 ;
        RECT 120.225 151.300 121.325 153.325 ;
        RECT 121.900 151.300 123.000 153.325 ;
        RECT 123.550 151.300 124.650 153.325 ;
        RECT 125.220 151.300 126.325 153.325 ;
        RECT 126.875 151.300 127.975 153.325 ;
        RECT 128.525 151.300 129.625 153.325 ;
        RECT 130.200 151.300 131.300 153.325 ;
        RECT 131.850 151.300 132.950 153.325 ;
        RECT 133.520 151.300 134.625 153.325 ;
        RECT 135.175 151.300 136.275 153.325 ;
        RECT 136.825 151.300 137.925 153.325 ;
        RECT 138.500 151.300 139.600 153.325 ;
        RECT 140.150 151.300 141.250 153.325 ;
        RECT 141.820 151.300 142.925 153.325 ;
        RECT 143.475 151.300 144.575 153.325 ;
        RECT 145.140 151.300 146.250 153.325 ;
        RECT 146.800 151.300 147.900 153.325 ;
        RECT 148.450 151.300 149.550 153.325 ;
        RECT 150.120 151.300 151.225 153.325 ;
        RECT 151.775 151.300 152.875 153.325 ;
        RECT 153.440 151.300 154.550 153.325 ;
        RECT 155.100 151.300 156.200 153.325 ;
        RECT 156.750 151.300 157.850 153.325 ;
        RECT 158.420 151.300 159.525 153.325 ;
        RECT 160.075 151.300 161.175 153.325 ;
        RECT 161.725 151.300 162.825 153.325 ;
        RECT 163.400 151.300 164.500 153.325 ;
        RECT 165.050 151.300 166.150 153.325 ;
        RECT 166.720 151.300 167.825 153.325 ;
        RECT 168.375 151.300 169.475 153.325 ;
        RECT 170.025 151.300 171.125 153.325 ;
        RECT 171.675 151.300 172.780 153.325 ;
        RECT 173.350 151.300 174.450 153.325 ;
        RECT 175.020 151.300 176.125 153.325 ;
        RECT 176.675 151.300 177.775 153.325 ;
        RECT 178.325 151.300 179.425 153.325 ;
        RECT 113.600 151.260 113.850 151.300 ;
        RECT 114.430 151.260 114.680 151.300 ;
        RECT 115.260 151.260 115.510 151.300 ;
        RECT 116.090 151.260 116.340 151.300 ;
        RECT 116.920 151.260 117.170 151.300 ;
        RECT 117.750 151.260 118.000 151.300 ;
        RECT 118.580 151.260 118.830 151.300 ;
        RECT 119.410 151.260 119.660 151.300 ;
        RECT 120.240 151.260 120.490 151.300 ;
        RECT 121.070 151.260 121.320 151.300 ;
        RECT 121.900 151.260 122.150 151.300 ;
        RECT 122.730 151.260 122.980 151.300 ;
        RECT 123.560 151.260 123.810 151.300 ;
        RECT 124.390 151.260 124.640 151.300 ;
        RECT 125.220 151.260 125.470 151.300 ;
        RECT 126.050 151.260 126.300 151.300 ;
        RECT 126.880 151.260 127.130 151.300 ;
        RECT 127.710 151.260 127.960 151.300 ;
        RECT 128.540 151.260 128.790 151.300 ;
        RECT 129.370 151.260 129.620 151.300 ;
        RECT 130.200 151.260 130.450 151.300 ;
        RECT 131.030 151.260 131.280 151.300 ;
        RECT 131.860 151.260 132.110 151.300 ;
        RECT 132.690 151.260 132.940 151.300 ;
        RECT 133.520 151.260 133.770 151.300 ;
        RECT 134.350 151.260 134.600 151.300 ;
        RECT 135.180 151.260 135.430 151.300 ;
        RECT 136.010 151.260 136.260 151.300 ;
        RECT 136.840 151.260 137.090 151.300 ;
        RECT 137.670 151.260 137.920 151.300 ;
        RECT 138.500 151.260 138.750 151.300 ;
        RECT 139.330 151.260 139.580 151.300 ;
        RECT 140.160 151.260 140.410 151.300 ;
        RECT 140.990 151.260 141.240 151.300 ;
        RECT 141.820 151.260 142.070 151.300 ;
        RECT 142.650 151.260 142.900 151.300 ;
        RECT 143.480 151.260 143.730 151.300 ;
        RECT 144.310 151.260 144.560 151.300 ;
        RECT 145.140 151.260 145.390 151.300 ;
        RECT 145.970 151.260 146.220 151.300 ;
        RECT 146.800 151.260 147.050 151.300 ;
        RECT 147.630 151.260 147.880 151.300 ;
        RECT 148.460 151.260 148.710 151.300 ;
        RECT 149.290 151.260 149.540 151.300 ;
        RECT 150.120 151.260 150.370 151.300 ;
        RECT 150.950 151.260 151.200 151.300 ;
        RECT 151.780 151.260 152.030 151.300 ;
        RECT 152.610 151.260 152.860 151.300 ;
        RECT 153.440 151.260 153.690 151.300 ;
        RECT 154.270 151.260 154.520 151.300 ;
        RECT 155.100 151.260 155.350 151.300 ;
        RECT 155.930 151.260 156.180 151.300 ;
        RECT 156.760 151.260 157.010 151.300 ;
        RECT 157.590 151.260 157.840 151.300 ;
        RECT 158.420 151.260 158.670 151.300 ;
        RECT 159.250 151.260 159.500 151.300 ;
        RECT 160.080 151.260 160.330 151.300 ;
        RECT 160.910 151.260 161.160 151.300 ;
        RECT 161.740 151.260 161.990 151.300 ;
        RECT 162.570 151.260 162.820 151.300 ;
        RECT 163.400 151.260 163.650 151.300 ;
        RECT 164.230 151.260 164.480 151.300 ;
        RECT 165.060 151.260 165.310 151.300 ;
        RECT 165.890 151.260 166.140 151.300 ;
        RECT 166.720 151.260 166.970 151.300 ;
        RECT 167.550 151.260 167.800 151.300 ;
        RECT 168.380 151.260 168.630 151.300 ;
        RECT 169.210 151.260 169.460 151.300 ;
        RECT 170.040 151.260 170.290 151.300 ;
        RECT 170.870 151.260 171.120 151.300 ;
        RECT 171.700 151.260 171.950 151.300 ;
        RECT 172.530 151.260 172.780 151.300 ;
        RECT 173.360 151.260 173.610 151.300 ;
        RECT 174.190 151.260 174.440 151.300 ;
        RECT 175.020 151.260 175.270 151.300 ;
        RECT 175.850 151.260 176.100 151.300 ;
        RECT 176.680 151.260 176.930 151.300 ;
        RECT 177.510 151.260 177.760 151.300 ;
        RECT 178.340 151.260 178.590 151.300 ;
        RECT 179.170 151.260 179.420 151.300 ;
        RECT 179.900 151.250 180.350 153.375 ;
        RECT 180.650 151.250 181.250 153.375 ;
        RECT 181.660 153.325 181.910 153.365 ;
        RECT 182.490 153.325 182.740 153.365 ;
        RECT 183.320 153.325 183.570 153.365 ;
        RECT 184.150 153.325 184.400 153.365 ;
        RECT 184.980 153.325 185.230 153.365 ;
        RECT 185.810 153.325 186.060 153.365 ;
        RECT 186.640 153.325 186.890 153.365 ;
        RECT 187.470 153.325 187.720 153.365 ;
        RECT 188.300 153.325 188.550 153.365 ;
        RECT 189.130 153.325 189.380 153.365 ;
        RECT 189.960 153.325 190.210 153.365 ;
        RECT 190.790 153.325 191.040 153.365 ;
        RECT 191.620 153.325 191.870 153.365 ;
        RECT 192.450 153.325 192.700 153.365 ;
        RECT 193.280 153.325 193.530 153.365 ;
        RECT 194.110 153.325 194.360 153.365 ;
        RECT 194.940 153.325 195.190 153.365 ;
        RECT 195.770 153.325 196.020 153.365 ;
        RECT 196.600 153.325 196.850 153.365 ;
        RECT 197.430 153.325 197.680 153.365 ;
        RECT 198.260 153.325 198.510 153.365 ;
        RECT 199.090 153.325 199.340 153.365 ;
        RECT 199.920 153.325 200.170 153.365 ;
        RECT 200.750 153.325 201.000 153.365 ;
        RECT 201.580 153.325 201.830 153.365 ;
        RECT 202.410 153.325 202.660 153.365 ;
        RECT 203.240 153.325 203.490 153.365 ;
        RECT 204.070 153.325 204.320 153.365 ;
        RECT 204.900 153.325 205.150 153.365 ;
        RECT 205.730 153.325 205.980 153.365 ;
        RECT 206.560 153.325 206.810 153.365 ;
        RECT 207.390 153.325 207.640 153.365 ;
        RECT 208.220 153.325 208.470 153.365 ;
        RECT 209.050 153.325 209.300 153.365 ;
        RECT 209.880 153.325 210.130 153.365 ;
        RECT 210.710 153.325 210.960 153.365 ;
        RECT 211.540 153.325 211.790 153.365 ;
        RECT 181.650 151.300 182.750 153.325 ;
        RECT 183.320 151.300 184.425 153.325 ;
        RECT 184.975 151.300 186.075 153.325 ;
        RECT 186.640 151.300 187.750 153.325 ;
        RECT 188.300 151.300 189.400 153.325 ;
        RECT 189.950 151.300 191.050 153.325 ;
        RECT 191.600 151.300 192.700 153.325 ;
        RECT 193.275 151.300 194.375 153.325 ;
        RECT 194.925 151.300 196.025 153.325 ;
        RECT 196.575 151.300 197.680 153.325 ;
        RECT 198.250 151.300 199.350 153.325 ;
        RECT 199.920 151.300 201.025 153.325 ;
        RECT 201.575 151.300 202.675 153.325 ;
        RECT 203.225 151.300 204.325 153.325 ;
        RECT 204.900 151.300 206.000 153.325 ;
        RECT 206.550 151.300 207.650 153.325 ;
        RECT 208.200 151.300 209.300 153.325 ;
        RECT 209.875 151.300 210.975 153.325 ;
        RECT 211.525 151.300 214.125 153.325 ;
        RECT 181.660 151.260 181.910 151.300 ;
        RECT 182.490 151.260 182.740 151.300 ;
        RECT 183.320 151.260 183.570 151.300 ;
        RECT 184.150 151.260 184.400 151.300 ;
        RECT 184.980 151.260 185.230 151.300 ;
        RECT 185.810 151.260 186.060 151.300 ;
        RECT 186.640 151.260 186.890 151.300 ;
        RECT 187.470 151.260 187.720 151.300 ;
        RECT 188.300 151.260 188.550 151.300 ;
        RECT 189.130 151.260 189.380 151.300 ;
        RECT 189.960 151.260 190.210 151.300 ;
        RECT 190.790 151.260 191.040 151.300 ;
        RECT 191.620 151.260 191.870 151.300 ;
        RECT 192.450 151.260 192.700 151.300 ;
        RECT 193.280 151.260 193.530 151.300 ;
        RECT 194.110 151.260 194.360 151.300 ;
        RECT 194.940 151.260 195.190 151.300 ;
        RECT 195.770 151.260 196.020 151.300 ;
        RECT 196.600 151.260 196.850 151.300 ;
        RECT 197.430 151.260 197.680 151.300 ;
        RECT 198.260 151.260 198.510 151.300 ;
        RECT 199.090 151.260 199.340 151.300 ;
        RECT 199.920 151.260 200.170 151.300 ;
        RECT 200.750 151.260 201.000 151.300 ;
        RECT 201.580 151.260 201.830 151.300 ;
        RECT 202.410 151.260 202.660 151.300 ;
        RECT 203.240 151.260 203.490 151.300 ;
        RECT 204.070 151.260 204.320 151.300 ;
        RECT 204.900 151.260 205.150 151.300 ;
        RECT 205.730 151.260 205.980 151.300 ;
        RECT 206.560 151.260 206.810 151.300 ;
        RECT 207.390 151.260 207.640 151.300 ;
        RECT 208.220 151.260 208.470 151.300 ;
        RECT 209.050 151.260 209.300 151.300 ;
        RECT 209.880 151.260 210.130 151.300 ;
        RECT 210.710 151.260 210.960 151.300 ;
        RECT 211.540 151.260 211.790 151.300 ;
        RECT 215.625 150.600 228.050 154.000 ;
        RECT 65.000 149.895 75.900 149.900 ;
        RECT 65.000 149.145 226.130 149.895 ;
        RECT 65.000 148.175 84.705 149.145 ;
        RECT 75.280 147.095 84.705 148.175 ;
        RECT 75.280 137.795 77.805 147.095 ;
        RECT 78.305 137.795 79.105 146.820 ;
        RECT 79.580 137.795 80.380 147.095 ;
        RECT 80.855 137.795 81.655 146.820 ;
        RECT 82.155 137.795 84.705 147.095 ;
        RECT 86.030 149.120 98.030 149.145 ;
        RECT 86.030 146.820 86.780 149.120 ;
        RECT 87.030 147.250 87.880 148.670 ;
        RECT 88.230 148.320 95.805 149.120 ;
        RECT 87.030 147.020 87.990 147.250 ;
        RECT 88.130 147.095 95.905 147.895 ;
        RECT 96.155 147.250 97.005 148.670 ;
        RECT 88.130 146.820 88.580 147.095 ;
        RECT 86.030 137.795 87.855 146.820 ;
        RECT 88.030 137.795 88.580 146.820 ;
        RECT 89.055 137.795 89.855 146.820 ;
        RECT 90.330 137.795 91.130 147.095 ;
        RECT 91.630 137.795 92.430 146.820 ;
        RECT 92.930 137.795 93.730 147.095 ;
        RECT 95.480 146.820 95.905 147.095 ;
        RECT 96.060 147.020 97.020 147.250 ;
        RECT 97.255 146.820 98.030 149.120 ;
        RECT 94.205 137.795 95.005 146.820 ;
        RECT 95.480 137.795 96.280 146.820 ;
        RECT 97.105 146.815 98.030 146.820 ;
        RECT 97.070 137.815 98.030 146.815 ;
        RECT 97.105 137.795 98.030 137.815 ;
        RECT 99.355 149.120 111.355 149.145 ;
        RECT 99.355 146.820 100.105 149.120 ;
        RECT 100.355 147.250 101.205 148.670 ;
        RECT 101.555 148.320 109.130 149.120 ;
        RECT 100.355 147.020 101.315 147.250 ;
        RECT 101.455 147.095 109.230 147.895 ;
        RECT 109.480 147.250 110.330 148.670 ;
        RECT 101.455 146.820 101.905 147.095 ;
        RECT 99.355 137.795 101.180 146.820 ;
        RECT 101.355 137.795 101.905 146.820 ;
        RECT 102.380 137.795 103.180 146.820 ;
        RECT 103.655 137.795 104.455 147.095 ;
        RECT 104.955 137.795 105.755 146.820 ;
        RECT 106.255 137.795 107.055 147.095 ;
        RECT 108.805 146.820 109.230 147.095 ;
        RECT 109.385 147.020 110.345 147.250 ;
        RECT 110.580 146.820 111.355 149.120 ;
        RECT 107.530 137.795 108.330 146.820 ;
        RECT 108.805 137.795 109.605 146.820 ;
        RECT 110.430 146.815 111.355 146.820 ;
        RECT 110.395 137.815 111.355 146.815 ;
        RECT 110.430 137.795 111.355 137.815 ;
        RECT 112.680 149.095 122.105 149.145 ;
        RECT 112.680 146.820 113.405 149.095 ;
        RECT 113.680 147.250 114.530 148.670 ;
        RECT 114.880 148.170 119.880 149.095 ;
        RECT 113.680 147.020 114.640 147.250 ;
        RECT 114.780 147.095 119.980 147.895 ;
        RECT 120.180 147.250 121.030 148.670 ;
        RECT 114.780 146.820 115.205 147.095 ;
        RECT 112.680 137.795 114.505 146.820 ;
        RECT 114.680 137.795 115.205 146.820 ;
        RECT 115.705 137.795 116.505 146.820 ;
        RECT 116.980 137.795 117.780 147.095 ;
        RECT 119.555 146.820 119.980 147.095 ;
        RECT 120.130 147.020 121.090 147.250 ;
        RECT 121.305 146.820 122.105 149.095 ;
        RECT 118.255 137.795 119.055 146.820 ;
        RECT 119.555 137.795 120.355 146.820 ;
        RECT 121.180 146.815 122.105 146.820 ;
        RECT 121.140 137.815 122.105 146.815 ;
        RECT 121.155 137.795 122.105 137.815 ;
        RECT 123.430 149.120 135.430 149.145 ;
        RECT 123.430 146.820 124.180 149.120 ;
        RECT 124.430 147.250 125.280 148.670 ;
        RECT 125.630 148.320 133.205 149.120 ;
        RECT 124.430 147.020 125.390 147.250 ;
        RECT 125.530 147.095 133.305 147.895 ;
        RECT 133.555 147.250 134.405 148.670 ;
        RECT 125.530 146.820 125.980 147.095 ;
        RECT 123.430 137.795 125.255 146.820 ;
        RECT 125.430 137.795 125.980 146.820 ;
        RECT 126.455 137.795 127.255 146.820 ;
        RECT 127.730 137.795 128.530 147.095 ;
        RECT 129.030 137.795 129.830 146.820 ;
        RECT 130.330 137.795 131.130 147.095 ;
        RECT 132.880 146.820 133.305 147.095 ;
        RECT 133.460 147.020 134.420 147.250 ;
        RECT 134.655 146.820 135.430 149.120 ;
        RECT 131.605 137.795 132.405 146.820 ;
        RECT 132.880 137.795 133.680 146.820 ;
        RECT 134.505 146.815 135.430 146.820 ;
        RECT 134.470 137.815 135.430 146.815 ;
        RECT 134.505 137.795 135.430 137.815 ;
        RECT 136.755 149.120 148.755 149.145 ;
        RECT 136.755 146.820 137.505 149.120 ;
        RECT 137.755 147.250 138.605 148.670 ;
        RECT 138.955 148.320 146.530 149.120 ;
        RECT 137.755 147.020 138.715 147.250 ;
        RECT 138.855 147.095 146.630 147.895 ;
        RECT 146.880 147.250 147.730 148.670 ;
        RECT 138.855 146.820 139.305 147.095 ;
        RECT 136.755 137.795 138.580 146.820 ;
        RECT 138.755 137.795 139.305 146.820 ;
        RECT 139.780 137.795 140.580 146.820 ;
        RECT 141.055 137.795 141.855 147.095 ;
        RECT 142.355 137.795 143.155 146.820 ;
        RECT 143.655 137.795 144.455 147.095 ;
        RECT 146.205 146.820 146.630 147.095 ;
        RECT 146.785 147.020 147.745 147.250 ;
        RECT 147.980 146.820 148.755 149.120 ;
        RECT 144.930 137.795 145.730 146.820 ;
        RECT 146.205 137.795 147.005 146.820 ;
        RECT 147.830 146.815 148.755 146.820 ;
        RECT 147.795 137.815 148.755 146.815 ;
        RECT 147.830 137.795 148.755 137.815 ;
        RECT 150.080 149.120 162.080 149.145 ;
        RECT 150.080 146.820 150.830 149.120 ;
        RECT 151.080 147.250 151.930 148.670 ;
        RECT 152.280 148.320 159.855 149.120 ;
        RECT 151.080 147.020 152.040 147.250 ;
        RECT 152.180 147.095 159.955 147.895 ;
        RECT 160.205 147.250 161.055 148.670 ;
        RECT 152.180 146.820 152.630 147.095 ;
        RECT 150.080 137.795 151.905 146.820 ;
        RECT 152.080 137.795 152.630 146.820 ;
        RECT 153.105 137.795 153.905 146.820 ;
        RECT 154.380 137.795 155.180 147.095 ;
        RECT 155.680 137.795 156.480 146.820 ;
        RECT 156.980 137.795 157.780 147.095 ;
        RECT 159.530 146.820 159.955 147.095 ;
        RECT 160.110 147.020 161.070 147.250 ;
        RECT 161.305 146.820 162.080 149.120 ;
        RECT 158.255 137.795 159.055 146.820 ;
        RECT 159.530 137.795 160.330 146.820 ;
        RECT 161.155 146.815 162.080 146.820 ;
        RECT 161.120 137.815 162.080 146.815 ;
        RECT 161.155 137.795 162.080 137.815 ;
        RECT 163.405 149.120 175.405 149.145 ;
        RECT 163.405 146.820 164.155 149.120 ;
        RECT 164.405 147.250 165.255 148.670 ;
        RECT 165.605 148.320 173.180 149.120 ;
        RECT 164.405 147.020 165.365 147.250 ;
        RECT 165.505 147.095 173.280 147.895 ;
        RECT 173.530 147.250 174.380 148.670 ;
        RECT 165.505 146.820 165.955 147.095 ;
        RECT 163.405 137.795 165.230 146.820 ;
        RECT 165.405 137.795 165.955 146.820 ;
        RECT 166.430 137.795 167.230 146.820 ;
        RECT 167.705 137.795 168.505 147.095 ;
        RECT 169.005 137.795 169.805 146.820 ;
        RECT 170.305 137.795 171.105 147.095 ;
        RECT 172.855 146.820 173.280 147.095 ;
        RECT 173.435 147.020 174.395 147.250 ;
        RECT 174.630 146.820 175.405 149.120 ;
        RECT 171.580 137.795 172.380 146.820 ;
        RECT 172.855 137.795 173.655 146.820 ;
        RECT 174.480 146.815 175.405 146.820 ;
        RECT 174.445 137.815 175.405 146.815 ;
        RECT 174.480 137.795 175.405 137.815 ;
        RECT 176.730 149.120 188.730 149.145 ;
        RECT 176.730 146.820 177.480 149.120 ;
        RECT 177.730 147.250 178.580 148.670 ;
        RECT 178.930 148.320 186.505 149.120 ;
        RECT 177.730 147.020 178.690 147.250 ;
        RECT 178.830 147.095 186.605 147.895 ;
        RECT 186.855 147.250 187.705 148.670 ;
        RECT 178.830 146.820 179.280 147.095 ;
        RECT 176.730 137.795 178.555 146.820 ;
        RECT 178.730 137.795 179.280 146.820 ;
        RECT 179.755 137.795 180.555 146.820 ;
        RECT 181.030 137.795 181.830 147.095 ;
        RECT 182.330 137.795 183.130 146.820 ;
        RECT 183.630 137.795 184.430 147.095 ;
        RECT 186.180 146.820 186.605 147.095 ;
        RECT 186.760 147.020 187.720 147.250 ;
        RECT 187.955 146.820 188.730 149.120 ;
        RECT 184.905 137.795 185.705 146.820 ;
        RECT 186.180 137.795 186.980 146.820 ;
        RECT 187.805 146.815 188.730 146.820 ;
        RECT 187.770 137.815 188.730 146.815 ;
        RECT 187.805 137.795 188.730 137.815 ;
        RECT 190.055 149.095 199.480 149.145 ;
        RECT 190.055 146.820 190.780 149.095 ;
        RECT 191.055 147.250 191.905 148.670 ;
        RECT 192.255 148.170 197.255 149.095 ;
        RECT 191.055 147.020 192.015 147.250 ;
        RECT 192.155 147.095 197.355 147.895 ;
        RECT 197.555 147.250 198.405 148.670 ;
        RECT 192.155 146.820 192.580 147.095 ;
        RECT 190.055 137.795 191.880 146.820 ;
        RECT 192.055 137.795 192.580 146.820 ;
        RECT 193.080 137.795 193.880 146.820 ;
        RECT 194.355 137.795 195.155 147.095 ;
        RECT 196.930 146.820 197.355 147.095 ;
        RECT 197.505 147.020 198.465 147.250 ;
        RECT 198.680 146.820 199.480 149.095 ;
        RECT 195.630 137.795 196.430 146.820 ;
        RECT 196.930 137.795 197.730 146.820 ;
        RECT 198.555 146.815 199.480 146.820 ;
        RECT 198.515 137.815 199.480 146.815 ;
        RECT 198.530 137.795 199.480 137.815 ;
        RECT 200.805 149.120 212.805 149.145 ;
        RECT 200.805 146.820 201.555 149.120 ;
        RECT 201.805 147.250 202.655 148.670 ;
        RECT 203.005 148.320 210.580 149.120 ;
        RECT 201.805 147.020 202.765 147.250 ;
        RECT 202.905 147.095 210.680 147.895 ;
        RECT 210.930 147.250 211.780 148.670 ;
        RECT 202.905 146.820 203.355 147.095 ;
        RECT 200.805 137.795 202.630 146.820 ;
        RECT 202.805 137.795 203.355 146.820 ;
        RECT 203.830 137.795 204.630 146.820 ;
        RECT 205.105 137.795 205.905 147.095 ;
        RECT 206.405 137.795 207.205 146.820 ;
        RECT 207.705 137.795 208.505 147.095 ;
        RECT 210.255 146.820 210.680 147.095 ;
        RECT 210.835 147.020 211.795 147.250 ;
        RECT 212.030 146.820 212.805 149.120 ;
        RECT 208.980 137.795 209.780 146.820 ;
        RECT 210.255 137.795 211.055 146.820 ;
        RECT 211.880 146.815 212.805 146.820 ;
        RECT 211.845 137.815 212.805 146.815 ;
        RECT 211.880 137.795 212.805 137.815 ;
        RECT 214.130 149.120 226.130 149.145 ;
        RECT 214.130 146.820 214.880 149.120 ;
        RECT 215.130 147.250 215.980 148.670 ;
        RECT 216.330 148.320 223.905 149.120 ;
        RECT 215.130 147.020 216.090 147.250 ;
        RECT 216.230 147.095 224.005 147.895 ;
        RECT 224.255 147.250 225.105 148.670 ;
        RECT 216.230 146.820 216.680 147.095 ;
        RECT 214.130 137.795 215.955 146.820 ;
        RECT 216.130 137.795 216.680 146.820 ;
        RECT 217.155 137.795 217.955 146.820 ;
        RECT 218.430 137.795 219.230 147.095 ;
        RECT 219.730 137.795 220.530 146.820 ;
        RECT 221.030 137.795 221.830 147.095 ;
        RECT 223.580 146.820 224.005 147.095 ;
        RECT 224.160 147.020 225.120 147.250 ;
        RECT 225.355 146.820 226.130 149.120 ;
        RECT 222.305 137.795 223.105 146.820 ;
        RECT 223.580 137.795 224.380 146.820 ;
        RECT 225.205 146.815 226.130 146.820 ;
        RECT 225.170 137.815 226.130 146.815 ;
        RECT 225.205 137.795 226.130 137.815 ;
        RECT 226.800 143.200 228.050 150.600 ;
        RECT 228.675 143.650 229.275 161.075 ;
        RECT 230.000 153.975 230.600 207.300 ;
        RECT 233.250 167.050 233.850 210.575 ;
        RECT 236.500 170.300 237.100 213.850 ;
        RECT 236.500 169.700 276.375 170.300 ;
        RECT 233.250 166.450 273.400 167.050 ;
        RECT 240.650 159.850 243.525 160.000 ;
        RECT 231.050 158.995 266.400 159.850 ;
        RECT 231.045 158.650 266.400 158.995 ;
        RECT 231.045 158.645 234.650 158.650 ;
        RECT 235.645 158.645 248.450 158.650 ;
        RECT 231.050 158.625 234.650 158.645 ;
        RECT 231.050 157.900 232.050 158.625 ;
        RECT 233.650 158.445 234.650 158.625 ;
        RECT 233.645 158.120 234.650 158.445 ;
        RECT 233.650 157.900 234.650 158.120 ;
        RECT 231.050 157.895 232.275 157.900 ;
        RECT 231.050 154.900 232.480 157.895 ;
        RECT 232.675 154.900 233.025 157.900 ;
        RECT 233.425 157.895 234.650 157.900 ;
        RECT 233.210 154.900 234.650 157.895 ;
        RECT 235.650 158.625 248.450 158.645 ;
        RECT 235.650 157.900 236.650 158.625 ;
        RECT 238.250 158.445 241.525 158.625 ;
        RECT 242.575 158.445 245.850 158.625 ;
        RECT 247.450 158.445 248.450 158.625 ;
        RECT 238.245 158.125 241.525 158.445 ;
        RECT 238.245 158.120 241.250 158.125 ;
        RECT 242.570 158.120 245.850 158.445 ;
        RECT 247.445 158.120 248.450 158.445 ;
        RECT 238.250 157.900 241.250 158.120 ;
        RECT 242.850 157.900 245.850 158.120 ;
        RECT 247.450 157.900 248.450 158.120 ;
        RECT 235.650 157.895 236.875 157.900 ;
        RECT 235.650 154.900 237.080 157.895 ;
        RECT 237.275 154.900 237.625 157.900 ;
        RECT 238.025 157.895 241.475 157.900 ;
        RECT 237.810 154.900 241.680 157.895 ;
        RECT 241.875 154.900 242.225 157.900 ;
        RECT 242.625 157.895 246.075 157.900 ;
        RECT 242.410 154.900 246.280 157.895 ;
        RECT 246.475 154.900 246.825 157.900 ;
        RECT 247.225 157.895 248.450 157.900 ;
        RECT 247.010 154.900 248.450 157.895 ;
        RECT 249.450 158.450 250.450 158.650 ;
        RECT 249.450 158.125 250.455 158.450 ;
        RECT 249.450 157.900 250.450 158.125 ;
        RECT 249.450 154.900 250.880 157.900 ;
        RECT 251.075 154.900 251.400 157.900 ;
        RECT 251.600 154.900 251.850 158.650 ;
        RECT 252.050 154.900 252.375 157.900 ;
        RECT 252.550 154.900 252.800 158.650 ;
        RECT 253.950 158.500 266.400 158.650 ;
        RECT 253.950 157.900 254.950 158.500 ;
        RECT 253.000 154.900 253.325 157.900 ;
        RECT 253.530 154.900 254.950 157.900 ;
        RECT 231.770 154.895 232.000 154.900 ;
        RECT 232.250 154.895 232.480 154.900 ;
        RECT 232.730 154.895 232.960 154.900 ;
        RECT 233.210 154.895 233.440 154.900 ;
        RECT 233.690 154.895 233.920 154.900 ;
        RECT 236.370 154.895 236.600 154.900 ;
        RECT 236.850 154.895 237.080 154.900 ;
        RECT 237.330 154.895 237.560 154.900 ;
        RECT 237.810 154.895 238.040 154.900 ;
        RECT 238.290 154.895 238.520 154.900 ;
        RECT 240.970 154.895 241.200 154.900 ;
        RECT 241.450 154.895 241.680 154.900 ;
        RECT 241.930 154.895 242.160 154.900 ;
        RECT 242.410 154.895 242.640 154.900 ;
        RECT 242.890 154.895 243.120 154.900 ;
        RECT 245.570 154.895 245.800 154.900 ;
        RECT 246.050 154.895 246.280 154.900 ;
        RECT 246.530 154.895 246.760 154.900 ;
        RECT 247.010 154.895 247.240 154.900 ;
        RECT 247.490 154.895 247.720 154.900 ;
        RECT 232.450 154.695 233.250 154.700 ;
        RECT 237.050 154.695 237.850 154.700 ;
        RECT 242.100 154.695 242.475 154.700 ;
        RECT 246.250 154.695 247.050 154.700 ;
        RECT 232.445 154.320 233.250 154.695 ;
        RECT 237.045 154.320 237.850 154.695 ;
        RECT 242.095 154.320 242.475 154.695 ;
        RECT 246.245 154.320 247.050 154.695 ;
        RECT 232.450 153.975 233.250 154.320 ;
        RECT 237.050 153.975 237.850 154.320 ;
        RECT 242.100 153.975 242.475 154.320 ;
        RECT 246.250 153.975 247.050 154.320 ;
        RECT 250.825 154.325 253.580 154.700 ;
        RECT 250.825 153.975 253.575 154.325 ;
        RECT 230.000 153.375 233.250 153.975 ;
        RECT 234.900 153.375 237.850 153.975 ;
        RECT 239.500 153.375 242.475 153.975 ;
        RECT 244.775 153.375 247.050 153.975 ;
        RECT 248.700 153.375 253.575 153.975 ;
        RECT 230.000 144.675 230.600 153.375 ;
        RECT 232.450 152.700 233.250 153.375 ;
        RECT 237.050 152.700 237.850 153.375 ;
        RECT 242.100 152.700 242.475 153.375 ;
        RECT 246.250 152.700 247.050 153.375 ;
        RECT 250.825 153.025 253.575 153.375 ;
        RECT 250.825 152.700 253.580 153.025 ;
        RECT 256.625 152.950 271.250 153.300 ;
        RECT 231.050 151.500 232.485 152.500 ;
        RECT 232.675 151.500 233.025 152.500 ;
        RECT 233.215 151.500 237.085 152.500 ;
        RECT 237.275 151.500 237.625 152.500 ;
        RECT 237.815 151.500 239.250 152.500 ;
        RECT 231.050 150.800 232.050 151.500 ;
        RECT 233.650 150.800 236.650 151.500 ;
        RECT 238.250 150.800 239.250 151.500 ;
        RECT 240.250 151.500 241.685 152.500 ;
        RECT 241.875 151.500 242.225 152.500 ;
        RECT 242.415 151.500 243.850 152.500 ;
        RECT 240.250 151.300 241.250 151.500 ;
        RECT 242.850 151.300 243.850 151.500 ;
        RECT 240.250 150.800 241.525 151.300 ;
        RECT 242.575 150.800 243.850 151.300 ;
        RECT 244.850 151.500 246.285 152.500 ;
        RECT 246.475 151.500 246.825 152.500 ;
        RECT 247.015 151.500 250.880 152.500 ;
        RECT 251.075 151.500 251.400 152.500 ;
        RECT 244.850 150.800 245.850 151.500 ;
        RECT 247.450 151.475 250.880 151.500 ;
        RECT 247.450 150.800 250.875 151.475 ;
        RECT 251.600 150.800 251.850 152.500 ;
        RECT 252.050 151.500 252.375 152.500 ;
        RECT 252.550 150.800 252.800 152.500 ;
        RECT 253.000 151.500 253.325 152.500 ;
        RECT 253.525 150.800 254.950 152.500 ;
        RECT 256.625 152.400 271.250 152.775 ;
        RECT 231.050 150.450 254.955 150.800 ;
        RECT 231.050 149.700 233.700 149.705 ;
        RECT 231.050 149.350 254.955 149.700 ;
        RECT 231.050 145.600 231.425 149.350 ;
        RECT 231.950 148.800 232.800 149.180 ;
        RECT 231.775 144.675 232.025 148.625 ;
        RECT 232.200 145.600 232.550 148.625 ;
        RECT 232.725 144.675 232.975 148.625 ;
        RECT 233.325 145.600 233.700 149.350 ;
        RECT 235.645 149.345 248.450 149.350 ;
        RECT 235.650 149.325 248.450 149.345 ;
        RECT 235.650 148.600 236.650 149.325 ;
        RECT 238.250 149.145 241.525 149.325 ;
        RECT 242.575 149.145 245.850 149.325 ;
        RECT 247.450 149.145 248.450 149.325 ;
        RECT 238.245 148.825 241.525 149.145 ;
        RECT 238.245 148.820 241.250 148.825 ;
        RECT 242.570 148.820 245.850 149.145 ;
        RECT 247.445 148.820 248.450 149.145 ;
        RECT 238.250 148.600 241.250 148.820 ;
        RECT 242.850 148.600 245.850 148.820 ;
        RECT 247.450 148.600 248.450 148.820 ;
        RECT 235.650 148.595 236.875 148.600 ;
        RECT 235.650 145.600 237.080 148.595 ;
        RECT 237.275 145.600 237.625 148.600 ;
        RECT 238.025 148.595 241.475 148.600 ;
        RECT 237.810 145.600 241.680 148.595 ;
        RECT 241.875 145.600 242.225 148.600 ;
        RECT 242.625 148.595 246.075 148.600 ;
        RECT 242.410 145.600 246.280 148.595 ;
        RECT 246.475 145.600 246.825 148.600 ;
        RECT 247.225 148.595 248.450 148.600 ;
        RECT 247.010 145.600 248.450 148.595 ;
        RECT 249.450 149.150 250.450 149.350 ;
        RECT 249.450 148.825 250.455 149.150 ;
        RECT 249.450 148.600 250.450 148.825 ;
        RECT 249.450 145.600 250.880 148.600 ;
        RECT 251.075 145.600 251.400 148.600 ;
        RECT 251.600 145.600 251.850 149.350 ;
        RECT 252.050 145.600 252.375 148.600 ;
        RECT 252.550 145.600 252.800 149.350 ;
        RECT 253.950 148.600 254.950 149.350 ;
        RECT 253.000 145.600 253.325 148.600 ;
        RECT 253.530 145.600 254.950 148.600 ;
        RECT 256.625 145.600 256.975 152.400 ;
        RECT 257.540 152.395 259.290 152.400 ;
        RECT 268.590 152.395 270.340 152.400 ;
        RECT 257.345 152.125 257.575 152.195 ;
        RECT 257.825 152.125 258.055 152.195 ;
        RECT 258.305 152.125 258.535 152.195 ;
        RECT 258.785 152.125 259.015 152.195 ;
        RECT 259.265 152.125 259.495 152.195 ;
        RECT 259.745 152.125 259.975 152.195 ;
        RECT 257.300 150.950 259.500 152.125 ;
        RECT 259.700 150.950 260.025 152.125 ;
        RECT 257.345 149.195 257.575 150.950 ;
        RECT 257.825 149.195 258.055 150.950 ;
        RECT 258.305 149.195 258.535 150.950 ;
        RECT 258.785 149.195 259.015 150.950 ;
        RECT 259.225 150.925 259.500 150.950 ;
        RECT 259.225 149.200 259.550 150.925 ;
        RECT 259.265 149.195 259.495 149.200 ;
        RECT 259.745 149.195 259.975 150.950 ;
        RECT 260.225 150.375 260.455 152.195 ;
        RECT 260.705 152.125 260.935 152.195 ;
        RECT 260.650 150.950 260.975 152.125 ;
        RECT 260.175 149.200 260.500 150.375 ;
        RECT 260.225 149.195 260.455 149.200 ;
        RECT 260.705 149.195 260.935 150.950 ;
        RECT 261.185 150.375 261.415 152.195 ;
        RECT 261.665 152.125 261.895 152.195 ;
        RECT 261.625 150.950 261.950 152.125 ;
        RECT 261.125 149.200 261.475 150.375 ;
        RECT 261.185 149.195 261.415 149.200 ;
        RECT 261.665 149.195 261.895 150.950 ;
        RECT 262.145 150.375 262.375 152.195 ;
        RECT 262.625 152.125 262.855 152.195 ;
        RECT 262.575 150.950 262.900 152.125 ;
        RECT 262.100 149.200 262.425 150.375 ;
        RECT 262.145 149.195 262.375 149.200 ;
        RECT 262.625 149.195 262.855 150.950 ;
        RECT 263.105 150.375 263.335 152.195 ;
        RECT 263.585 152.125 263.815 152.195 ;
        RECT 263.525 150.950 263.875 152.125 ;
        RECT 263.050 149.200 263.375 150.375 ;
        RECT 263.105 149.195 263.335 149.200 ;
        RECT 263.585 149.195 263.815 150.950 ;
        RECT 264.065 150.375 264.295 152.195 ;
        RECT 264.545 152.125 264.775 152.195 ;
        RECT 264.500 150.950 264.825 152.125 ;
        RECT 264.025 149.200 264.350 150.375 ;
        RECT 264.065 149.195 264.295 149.200 ;
        RECT 264.545 149.195 264.775 150.950 ;
        RECT 265.025 150.375 265.255 152.195 ;
        RECT 265.505 152.125 265.735 152.195 ;
        RECT 265.450 150.950 265.775 152.125 ;
        RECT 264.975 149.200 265.300 150.375 ;
        RECT 265.025 149.195 265.255 149.200 ;
        RECT 265.505 149.195 265.735 150.950 ;
        RECT 265.985 150.375 266.215 152.195 ;
        RECT 266.465 152.125 266.695 152.195 ;
        RECT 266.425 150.950 266.750 152.125 ;
        RECT 265.925 149.200 266.250 150.375 ;
        RECT 265.985 149.195 266.215 149.200 ;
        RECT 266.465 149.195 266.695 150.950 ;
        RECT 266.945 150.375 267.175 152.195 ;
        RECT 267.425 152.125 267.655 152.195 ;
        RECT 267.375 150.950 267.700 152.125 ;
        RECT 266.900 149.200 267.225 150.375 ;
        RECT 266.945 149.195 267.175 149.200 ;
        RECT 267.425 149.195 267.655 150.950 ;
        RECT 267.905 150.375 268.135 152.195 ;
        RECT 268.385 152.125 268.615 152.195 ;
        RECT 268.865 152.125 269.095 152.195 ;
        RECT 269.345 152.125 269.575 152.195 ;
        RECT 269.825 152.125 270.055 152.195 ;
        RECT 270.305 152.125 270.535 152.195 ;
        RECT 268.325 150.950 270.575 152.125 ;
        RECT 267.850 149.200 268.175 150.375 ;
        RECT 267.905 149.195 268.135 149.200 ;
        RECT 268.385 149.195 268.615 150.950 ;
        RECT 268.865 149.195 269.095 150.950 ;
        RECT 269.345 149.195 269.575 150.950 ;
        RECT 269.825 149.195 270.055 150.950 ;
        RECT 270.305 149.195 270.535 150.950 ;
        RECT 257.525 147.000 270.350 149.000 ;
        RECT 257.345 146.150 257.575 146.800 ;
        RECT 257.825 146.150 258.055 146.800 ;
        RECT 258.305 146.150 258.535 146.800 ;
        RECT 258.785 146.150 259.015 146.800 ;
        RECT 259.225 146.175 259.550 146.800 ;
        RECT 259.225 146.150 259.525 146.175 ;
        RECT 259.745 146.150 259.975 146.800 ;
        RECT 260.175 146.400 260.500 146.800 ;
        RECT 257.300 145.750 259.525 146.150 ;
        RECT 259.700 145.750 260.025 146.150 ;
        RECT 260.225 145.800 260.455 146.400 ;
        RECT 260.705 146.150 260.935 146.800 ;
        RECT 261.125 146.400 261.475 146.800 ;
        RECT 260.650 145.750 261.000 146.150 ;
        RECT 261.185 145.800 261.415 146.400 ;
        RECT 261.665 146.150 261.895 146.800 ;
        RECT 262.100 146.400 262.425 146.800 ;
        RECT 261.625 145.750 261.950 146.150 ;
        RECT 262.145 145.800 262.375 146.400 ;
        RECT 262.625 146.150 262.855 146.800 ;
        RECT 263.050 146.400 263.375 146.800 ;
        RECT 262.575 145.750 262.900 146.150 ;
        RECT 263.105 145.800 263.335 146.400 ;
        RECT 263.585 146.150 263.815 146.800 ;
        RECT 264.025 146.400 264.350 146.800 ;
        RECT 263.525 145.750 263.875 146.150 ;
        RECT 264.065 145.800 264.295 146.400 ;
        RECT 264.545 146.150 264.775 146.800 ;
        RECT 264.975 146.400 265.300 146.800 ;
        RECT 264.500 145.750 264.825 146.150 ;
        RECT 265.025 145.800 265.255 146.400 ;
        RECT 265.505 146.150 265.735 146.800 ;
        RECT 265.925 146.400 266.275 146.800 ;
        RECT 265.450 145.750 265.800 146.150 ;
        RECT 265.985 145.800 266.215 146.400 ;
        RECT 266.465 146.150 266.695 146.800 ;
        RECT 266.900 146.400 267.225 146.800 ;
        RECT 266.425 145.750 266.750 146.150 ;
        RECT 266.945 145.800 267.175 146.400 ;
        RECT 267.425 146.150 267.655 146.800 ;
        RECT 267.850 146.400 268.200 146.800 ;
        RECT 267.375 145.750 267.700 146.150 ;
        RECT 267.905 145.800 268.135 146.400 ;
        RECT 268.385 146.150 268.615 146.800 ;
        RECT 268.865 146.150 269.095 146.800 ;
        RECT 269.345 146.150 269.575 146.800 ;
        RECT 269.825 146.150 270.055 146.800 ;
        RECT 270.305 146.150 270.535 146.800 ;
        RECT 268.325 145.750 270.575 146.150 ;
        RECT 270.900 145.600 271.250 152.400 ;
        RECT 236.370 145.595 236.600 145.600 ;
        RECT 236.850 145.595 237.080 145.600 ;
        RECT 237.330 145.595 237.560 145.600 ;
        RECT 237.810 145.595 238.040 145.600 ;
        RECT 238.290 145.595 238.520 145.600 ;
        RECT 240.970 145.595 241.200 145.600 ;
        RECT 241.450 145.595 241.680 145.600 ;
        RECT 241.930 145.595 242.160 145.600 ;
        RECT 242.410 145.595 242.640 145.600 ;
        RECT 242.890 145.595 243.120 145.600 ;
        RECT 245.570 145.595 245.800 145.600 ;
        RECT 246.050 145.595 246.280 145.600 ;
        RECT 246.530 145.595 246.760 145.600 ;
        RECT 247.010 145.595 247.240 145.600 ;
        RECT 247.490 145.595 247.720 145.600 ;
        RECT 237.050 145.395 237.850 145.400 ;
        RECT 242.100 145.395 242.475 145.400 ;
        RECT 246.250 145.395 247.050 145.400 ;
        RECT 230.000 144.075 232.975 144.675 ;
        RECT 226.800 141.500 231.425 143.200 ;
        RECT 231.775 142.200 232.025 144.075 ;
        RECT 232.200 142.200 232.550 143.200 ;
        RECT 232.725 142.200 232.975 144.075 ;
        RECT 233.325 143.200 233.700 145.350 ;
        RECT 237.045 145.020 237.850 145.395 ;
        RECT 242.095 145.020 242.475 145.395 ;
        RECT 246.245 145.020 247.050 145.395 ;
        RECT 237.050 144.675 237.850 145.020 ;
        RECT 242.100 144.675 242.475 145.020 ;
        RECT 246.250 144.675 247.050 145.020 ;
        RECT 250.825 145.025 253.580 145.400 ;
        RECT 256.625 145.275 271.250 145.600 ;
        RECT 250.825 144.675 253.575 145.025 ;
        RECT 256.625 144.750 271.250 145.100 ;
        RECT 234.900 144.075 237.850 144.675 ;
        RECT 239.500 144.075 242.475 144.675 ;
        RECT 244.775 144.075 247.050 144.675 ;
        RECT 248.700 144.075 253.575 144.675 ;
        RECT 237.050 143.400 237.850 144.075 ;
        RECT 242.100 143.400 242.475 144.075 ;
        RECT 246.250 143.400 247.050 144.075 ;
        RECT 250.825 143.725 253.575 144.075 ;
        RECT 250.825 143.400 253.580 143.725 ;
        RECT 233.325 142.200 237.085 143.200 ;
        RECT 237.275 142.200 237.625 143.200 ;
        RECT 237.815 142.200 239.250 143.200 ;
        RECT 231.950 141.675 232.800 142.000 ;
        RECT 233.325 141.500 236.650 142.200 ;
        RECT 238.250 141.500 239.250 142.200 ;
        RECT 240.250 142.200 241.685 143.200 ;
        RECT 241.875 142.200 242.225 143.200 ;
        RECT 242.415 142.200 243.850 143.200 ;
        RECT 240.250 142.000 241.250 142.200 ;
        RECT 242.850 142.000 243.850 142.200 ;
        RECT 240.250 141.500 241.525 142.000 ;
        RECT 242.575 141.500 243.850 142.000 ;
        RECT 244.850 142.200 246.285 143.200 ;
        RECT 246.475 142.200 246.825 143.200 ;
        RECT 247.015 142.200 250.880 143.200 ;
        RECT 251.075 142.200 251.400 143.200 ;
        RECT 244.850 141.500 245.850 142.200 ;
        RECT 247.450 142.175 250.880 142.200 ;
        RECT 247.450 141.500 250.875 142.175 ;
        RECT 251.600 141.500 251.850 143.200 ;
        RECT 252.050 142.200 252.375 143.200 ;
        RECT 252.550 141.500 252.800 143.200 ;
        RECT 253.000 142.200 253.325 143.200 ;
        RECT 253.525 141.650 254.950 143.200 ;
        RECT 253.525 141.500 261.450 141.650 ;
        RECT 226.800 140.300 261.450 141.500 ;
        RECT 77.570 137.570 78.530 137.610 ;
        RECT 78.860 137.570 79.820 137.610 ;
        RECT 80.150 137.570 81.110 137.610 ;
        RECT 81.440 137.570 82.400 137.610 ;
        RECT 88.320 137.570 89.280 137.610 ;
        RECT 89.610 137.595 90.570 137.610 ;
        RECT 90.900 137.595 91.860 137.610 ;
        RECT 89.610 137.570 91.860 137.595 ;
        RECT 92.190 137.570 93.150 137.610 ;
        RECT 93.480 137.570 94.440 137.610 ;
        RECT 94.770 137.570 95.730 137.610 ;
        RECT 77.570 137.395 82.430 137.570 ;
        RECT 88.320 137.395 95.730 137.570 ;
        RECT 101.645 137.570 102.605 137.610 ;
        RECT 102.935 137.595 103.895 137.610 ;
        RECT 104.225 137.595 105.185 137.610 ;
        RECT 102.935 137.570 105.185 137.595 ;
        RECT 105.515 137.570 106.475 137.610 ;
        RECT 106.805 137.570 107.765 137.610 ;
        RECT 108.095 137.570 109.055 137.610 ;
        RECT 101.645 137.395 109.055 137.570 ;
        RECT 114.970 137.570 115.930 137.610 ;
        RECT 116.260 137.570 117.220 137.610 ;
        RECT 117.550 137.570 118.510 137.610 ;
        RECT 118.840 137.570 119.800 137.610 ;
        RECT 125.720 137.570 126.680 137.610 ;
        RECT 127.010 137.595 127.970 137.610 ;
        RECT 128.300 137.595 129.260 137.610 ;
        RECT 127.010 137.570 129.260 137.595 ;
        RECT 129.590 137.570 130.550 137.610 ;
        RECT 130.880 137.570 131.840 137.610 ;
        RECT 132.170 137.570 133.130 137.610 ;
        RECT 114.970 137.545 119.830 137.570 ;
        RECT 114.970 137.395 120.805 137.545 ;
        RECT 125.720 137.395 133.130 137.570 ;
        RECT 139.045 137.570 140.005 137.610 ;
        RECT 140.335 137.595 141.295 137.610 ;
        RECT 141.625 137.595 142.585 137.610 ;
        RECT 140.335 137.570 142.585 137.595 ;
        RECT 142.915 137.570 143.875 137.610 ;
        RECT 144.205 137.570 145.165 137.610 ;
        RECT 145.495 137.570 146.455 137.610 ;
        RECT 139.045 137.395 146.455 137.570 ;
        RECT 152.370 137.570 153.330 137.610 ;
        RECT 153.660 137.595 154.620 137.610 ;
        RECT 154.950 137.595 155.910 137.610 ;
        RECT 153.660 137.570 155.910 137.595 ;
        RECT 156.240 137.570 157.200 137.610 ;
        RECT 157.530 137.570 158.490 137.610 ;
        RECT 158.820 137.570 159.780 137.610 ;
        RECT 152.370 137.395 159.780 137.570 ;
        RECT 165.695 137.570 166.655 137.610 ;
        RECT 166.985 137.595 167.945 137.610 ;
        RECT 168.275 137.595 169.235 137.610 ;
        RECT 166.985 137.570 169.235 137.595 ;
        RECT 169.565 137.570 170.525 137.610 ;
        RECT 170.855 137.570 171.815 137.610 ;
        RECT 172.145 137.570 173.105 137.610 ;
        RECT 165.695 137.395 173.105 137.570 ;
        RECT 179.020 137.570 179.980 137.610 ;
        RECT 180.310 137.595 181.270 137.610 ;
        RECT 181.600 137.595 182.560 137.610 ;
        RECT 180.310 137.570 182.560 137.595 ;
        RECT 182.890 137.570 183.850 137.610 ;
        RECT 184.180 137.570 185.140 137.610 ;
        RECT 185.470 137.570 186.430 137.610 ;
        RECT 179.020 137.395 186.430 137.570 ;
        RECT 192.345 137.570 193.305 137.610 ;
        RECT 193.635 137.570 194.595 137.610 ;
        RECT 194.925 137.570 195.885 137.610 ;
        RECT 196.215 137.570 197.175 137.610 ;
        RECT 203.095 137.570 204.055 137.610 ;
        RECT 204.385 137.595 205.345 137.610 ;
        RECT 205.675 137.595 206.635 137.610 ;
        RECT 204.385 137.570 206.635 137.595 ;
        RECT 206.965 137.570 207.925 137.610 ;
        RECT 208.255 137.570 209.215 137.610 ;
        RECT 209.545 137.570 210.505 137.610 ;
        RECT 192.345 137.395 198.180 137.570 ;
        RECT 203.095 137.395 210.505 137.570 ;
        RECT 216.420 137.570 217.380 137.610 ;
        RECT 217.710 137.595 218.670 137.610 ;
        RECT 219.000 137.595 219.960 137.610 ;
        RECT 217.710 137.570 219.960 137.595 ;
        RECT 220.290 137.570 221.250 137.610 ;
        RECT 221.580 137.570 222.540 137.610 ;
        RECT 222.870 137.570 223.830 137.610 ;
        RECT 216.420 137.395 223.830 137.570 ;
        RECT 72.650 137.245 75.275 137.250 ;
        RECT 77.555 137.245 82.430 137.395 ;
        RECT 72.650 136.000 82.430 137.245 ;
        RECT 75.105 135.995 82.430 136.000 ;
        RECT 77.555 135.845 82.430 135.995 ;
        RECT 85.680 135.845 95.730 137.395 ;
        RECT 99.005 135.845 109.055 137.395 ;
        RECT 110.755 135.845 120.805 137.395 ;
        RECT 123.080 135.845 133.130 137.395 ;
        RECT 136.405 135.845 146.455 137.395 ;
        RECT 149.730 135.845 159.780 137.395 ;
        RECT 163.055 135.845 173.105 137.395 ;
        RECT 176.380 135.845 186.430 137.395 ;
        RECT 189.705 135.845 198.180 137.395 ;
        RECT 200.455 135.845 210.505 137.395 ;
        RECT 213.780 135.845 223.830 137.395 ;
        RECT 77.570 135.670 82.430 135.845 ;
        RECT 88.320 135.670 95.730 135.845 ;
        RECT 77.570 135.630 78.530 135.670 ;
        RECT 78.860 135.630 79.820 135.670 ;
        RECT 80.150 135.630 81.110 135.670 ;
        RECT 81.440 135.630 82.400 135.670 ;
        RECT 88.320 135.630 89.280 135.670 ;
        RECT 89.610 135.645 91.860 135.670 ;
        RECT 89.610 135.630 90.570 135.645 ;
        RECT 90.900 135.630 91.860 135.645 ;
        RECT 92.190 135.630 93.150 135.670 ;
        RECT 93.480 135.630 94.440 135.670 ;
        RECT 94.770 135.630 95.730 135.670 ;
        RECT 101.645 135.670 109.055 135.845 ;
        RECT 101.645 135.630 102.605 135.670 ;
        RECT 102.935 135.645 105.185 135.670 ;
        RECT 102.935 135.630 103.895 135.645 ;
        RECT 104.225 135.630 105.185 135.645 ;
        RECT 105.515 135.630 106.475 135.670 ;
        RECT 106.805 135.630 107.765 135.670 ;
        RECT 108.095 135.630 109.055 135.670 ;
        RECT 114.970 135.670 120.805 135.845 ;
        RECT 125.720 135.670 133.130 135.845 ;
        RECT 114.970 135.630 115.930 135.670 ;
        RECT 116.260 135.630 117.220 135.670 ;
        RECT 117.550 135.630 118.510 135.670 ;
        RECT 118.840 135.630 119.800 135.670 ;
        RECT 125.720 135.630 126.680 135.670 ;
        RECT 127.010 135.645 129.260 135.670 ;
        RECT 127.010 135.630 127.970 135.645 ;
        RECT 128.300 135.630 129.260 135.645 ;
        RECT 129.590 135.630 130.550 135.670 ;
        RECT 130.880 135.630 131.840 135.670 ;
        RECT 132.170 135.630 133.130 135.670 ;
        RECT 139.045 135.670 146.455 135.845 ;
        RECT 139.045 135.630 140.005 135.670 ;
        RECT 140.335 135.645 142.585 135.670 ;
        RECT 140.335 135.630 141.295 135.645 ;
        RECT 141.625 135.630 142.585 135.645 ;
        RECT 142.915 135.630 143.875 135.670 ;
        RECT 144.205 135.630 145.165 135.670 ;
        RECT 145.495 135.630 146.455 135.670 ;
        RECT 152.370 135.670 159.780 135.845 ;
        RECT 152.370 135.630 153.330 135.670 ;
        RECT 153.660 135.645 155.910 135.670 ;
        RECT 153.660 135.630 154.620 135.645 ;
        RECT 154.950 135.630 155.910 135.645 ;
        RECT 156.240 135.630 157.200 135.670 ;
        RECT 157.530 135.630 158.490 135.670 ;
        RECT 158.820 135.630 159.780 135.670 ;
        RECT 165.695 135.670 173.105 135.845 ;
        RECT 165.695 135.630 166.655 135.670 ;
        RECT 166.985 135.645 169.235 135.670 ;
        RECT 166.985 135.630 167.945 135.645 ;
        RECT 168.275 135.630 169.235 135.645 ;
        RECT 169.565 135.630 170.525 135.670 ;
        RECT 170.855 135.630 171.815 135.670 ;
        RECT 172.145 135.630 173.105 135.670 ;
        RECT 179.020 135.670 186.430 135.845 ;
        RECT 179.020 135.630 179.980 135.670 ;
        RECT 180.310 135.645 182.560 135.670 ;
        RECT 180.310 135.630 181.270 135.645 ;
        RECT 181.600 135.630 182.560 135.645 ;
        RECT 182.890 135.630 183.850 135.670 ;
        RECT 184.180 135.630 185.140 135.670 ;
        RECT 185.470 135.630 186.430 135.670 ;
        RECT 192.345 135.670 198.180 135.845 ;
        RECT 203.095 135.670 210.505 135.845 ;
        RECT 192.345 135.630 193.305 135.670 ;
        RECT 193.635 135.630 194.595 135.670 ;
        RECT 194.925 135.630 195.885 135.670 ;
        RECT 196.215 135.630 197.175 135.670 ;
        RECT 203.095 135.630 204.055 135.670 ;
        RECT 204.385 135.645 206.635 135.670 ;
        RECT 204.385 135.630 205.345 135.645 ;
        RECT 205.675 135.630 206.635 135.645 ;
        RECT 206.965 135.630 207.925 135.670 ;
        RECT 208.255 135.630 209.215 135.670 ;
        RECT 209.545 135.630 210.505 135.670 ;
        RECT 216.420 135.670 223.830 135.845 ;
        RECT 216.420 135.630 217.380 135.670 ;
        RECT 217.710 135.645 219.960 135.670 ;
        RECT 217.710 135.630 218.670 135.645 ;
        RECT 219.000 135.630 219.960 135.645 ;
        RECT 220.290 135.630 221.250 135.670 ;
        RECT 221.580 135.630 222.540 135.670 ;
        RECT 222.870 135.630 223.830 135.670 ;
        RECT 226.800 135.500 228.050 140.300 ;
        RECT 226.125 135.495 228.050 135.500 ;
        RECT 75.280 135.425 77.830 135.470 ;
        RECT 75.275 132.525 77.830 135.425 ;
        RECT 75.280 132.195 77.830 132.525 ;
        RECT 78.305 132.470 79.105 135.470 ;
        RECT 79.580 132.195 80.380 135.470 ;
        RECT 80.855 132.470 81.655 135.470 ;
        RECT 82.130 132.195 84.705 135.470 ;
        RECT 75.280 131.125 84.705 132.195 ;
        RECT 75.025 130.195 84.705 131.125 ;
        RECT 86.030 132.470 86.980 135.495 ;
        RECT 97.105 135.470 98.030 135.495 ;
        RECT 87.755 132.470 88.555 135.470 ;
        RECT 89.055 132.470 89.855 135.470 ;
        RECT 86.030 132.445 86.955 132.470 ;
        RECT 86.030 130.220 86.780 132.445 ;
        RECT 87.030 132.080 87.990 132.310 ;
        RECT 88.130 132.195 88.555 132.470 ;
        RECT 90.330 132.195 91.130 135.470 ;
        RECT 91.630 132.470 92.430 135.470 ;
        RECT 92.905 132.195 93.705 135.470 ;
        RECT 94.205 132.470 95.005 135.470 ;
        RECT 95.480 132.470 96.280 135.470 ;
        RECT 97.070 132.470 98.030 135.470 ;
        RECT 95.480 132.195 95.905 132.470 ;
        RECT 87.030 130.670 87.880 132.080 ;
        RECT 88.130 131.395 95.905 132.195 ;
        RECT 96.060 132.080 97.020 132.310 ;
        RECT 88.230 130.220 95.805 131.020 ;
        RECT 96.155 130.670 97.005 132.080 ;
        RECT 97.255 130.220 98.030 132.470 ;
        RECT 86.030 130.195 98.030 130.220 ;
        RECT 99.355 132.470 100.305 135.495 ;
        RECT 110.430 135.470 111.355 135.495 ;
        RECT 101.080 132.470 101.880 135.470 ;
        RECT 102.380 132.470 103.180 135.470 ;
        RECT 99.355 132.445 100.280 132.470 ;
        RECT 99.355 130.220 100.105 132.445 ;
        RECT 100.355 132.080 101.315 132.310 ;
        RECT 101.455 132.195 101.880 132.470 ;
        RECT 103.655 132.195 104.455 135.470 ;
        RECT 104.955 132.470 105.755 135.470 ;
        RECT 106.230 132.195 107.030 135.470 ;
        RECT 107.530 132.470 108.330 135.470 ;
        RECT 108.805 132.470 109.605 135.470 ;
        RECT 110.395 132.470 111.355 135.470 ;
        RECT 108.805 132.195 109.230 132.470 ;
        RECT 100.355 130.670 101.205 132.080 ;
        RECT 101.455 131.395 109.230 132.195 ;
        RECT 109.385 132.080 110.345 132.310 ;
        RECT 101.555 130.220 109.130 131.020 ;
        RECT 109.480 130.670 110.330 132.080 ;
        RECT 110.580 130.220 111.355 132.470 ;
        RECT 99.355 130.195 111.355 130.220 ;
        RECT 112.680 132.445 113.630 135.470 ;
        RECT 114.405 132.470 115.205 135.470 ;
        RECT 115.705 132.470 116.505 135.470 ;
        RECT 112.680 130.195 113.405 132.445 ;
        RECT 113.680 132.080 114.640 132.310 ;
        RECT 114.780 132.195 115.205 132.470 ;
        RECT 116.980 132.195 117.780 135.470 ;
        RECT 118.255 132.470 119.055 135.470 ;
        RECT 119.555 132.470 120.355 135.470 ;
        RECT 121.140 132.470 122.105 135.470 ;
        RECT 119.555 132.195 119.980 132.470 ;
        RECT 121.155 132.445 122.105 132.470 ;
        RECT 113.680 130.670 114.530 132.080 ;
        RECT 114.780 131.395 119.980 132.195 ;
        RECT 120.130 132.080 121.090 132.310 ;
        RECT 114.880 130.195 119.880 131.120 ;
        RECT 120.180 130.670 121.030 132.080 ;
        RECT 121.305 130.195 122.105 132.445 ;
        RECT 123.430 132.470 124.380 135.495 ;
        RECT 134.505 135.470 135.430 135.495 ;
        RECT 125.155 132.470 125.955 135.470 ;
        RECT 126.455 132.470 127.255 135.470 ;
        RECT 123.430 132.445 124.355 132.470 ;
        RECT 123.430 130.220 124.180 132.445 ;
        RECT 124.430 132.080 125.390 132.310 ;
        RECT 125.530 132.195 125.955 132.470 ;
        RECT 127.730 132.195 128.530 135.470 ;
        RECT 129.030 132.470 129.830 135.470 ;
        RECT 130.305 132.195 131.105 135.470 ;
        RECT 131.605 132.470 132.405 135.470 ;
        RECT 132.880 132.470 133.680 135.470 ;
        RECT 134.470 132.470 135.430 135.470 ;
        RECT 132.880 132.195 133.305 132.470 ;
        RECT 124.430 130.670 125.280 132.080 ;
        RECT 125.530 131.395 133.305 132.195 ;
        RECT 133.460 132.080 134.420 132.310 ;
        RECT 125.630 130.220 133.205 131.020 ;
        RECT 133.555 130.670 134.405 132.080 ;
        RECT 134.655 130.220 135.430 132.470 ;
        RECT 123.430 130.195 135.430 130.220 ;
        RECT 136.755 132.470 137.705 135.495 ;
        RECT 147.830 135.470 148.755 135.495 ;
        RECT 138.480 132.470 139.280 135.470 ;
        RECT 139.780 132.470 140.580 135.470 ;
        RECT 136.755 132.445 137.680 132.470 ;
        RECT 136.755 130.220 137.505 132.445 ;
        RECT 137.755 132.080 138.715 132.310 ;
        RECT 138.855 132.195 139.280 132.470 ;
        RECT 141.055 132.195 141.855 135.470 ;
        RECT 142.355 132.470 143.155 135.470 ;
        RECT 143.630 132.195 144.430 135.470 ;
        RECT 144.930 132.470 145.730 135.470 ;
        RECT 146.205 132.470 147.005 135.470 ;
        RECT 147.795 132.470 148.755 135.470 ;
        RECT 146.205 132.195 146.630 132.470 ;
        RECT 137.755 130.670 138.605 132.080 ;
        RECT 138.855 131.395 146.630 132.195 ;
        RECT 146.785 132.080 147.745 132.310 ;
        RECT 138.955 130.220 146.530 131.020 ;
        RECT 146.880 130.670 147.730 132.080 ;
        RECT 147.980 130.220 148.755 132.470 ;
        RECT 136.755 130.195 148.755 130.220 ;
        RECT 150.080 132.470 151.030 135.495 ;
        RECT 161.155 135.470 162.080 135.495 ;
        RECT 151.805 132.470 152.605 135.470 ;
        RECT 153.105 132.470 153.905 135.470 ;
        RECT 150.080 132.445 151.005 132.470 ;
        RECT 150.080 130.220 150.830 132.445 ;
        RECT 151.080 132.080 152.040 132.310 ;
        RECT 152.180 132.195 152.605 132.470 ;
        RECT 154.380 132.195 155.180 135.470 ;
        RECT 155.680 132.470 156.480 135.470 ;
        RECT 156.955 132.195 157.755 135.470 ;
        RECT 158.255 132.470 159.055 135.470 ;
        RECT 159.530 132.470 160.330 135.470 ;
        RECT 161.120 132.470 162.080 135.470 ;
        RECT 159.530 132.195 159.955 132.470 ;
        RECT 151.080 130.670 151.930 132.080 ;
        RECT 152.180 131.395 159.955 132.195 ;
        RECT 160.110 132.080 161.070 132.310 ;
        RECT 152.280 130.220 159.855 131.020 ;
        RECT 160.205 130.670 161.055 132.080 ;
        RECT 161.305 130.220 162.080 132.470 ;
        RECT 150.080 130.195 162.080 130.220 ;
        RECT 163.405 132.470 164.355 135.495 ;
        RECT 174.480 135.470 175.405 135.495 ;
        RECT 165.130 132.470 165.930 135.470 ;
        RECT 166.430 132.470 167.230 135.470 ;
        RECT 163.405 132.445 164.330 132.470 ;
        RECT 163.405 130.220 164.155 132.445 ;
        RECT 164.405 132.080 165.365 132.310 ;
        RECT 165.505 132.195 165.930 132.470 ;
        RECT 167.705 132.195 168.505 135.470 ;
        RECT 169.005 132.470 169.805 135.470 ;
        RECT 170.280 132.195 171.080 135.470 ;
        RECT 171.580 132.470 172.380 135.470 ;
        RECT 172.855 132.470 173.655 135.470 ;
        RECT 174.445 132.470 175.405 135.470 ;
        RECT 172.855 132.195 173.280 132.470 ;
        RECT 164.405 130.670 165.255 132.080 ;
        RECT 165.505 131.395 173.280 132.195 ;
        RECT 173.435 132.080 174.395 132.310 ;
        RECT 165.605 130.220 173.180 131.020 ;
        RECT 173.530 130.670 174.380 132.080 ;
        RECT 174.630 130.220 175.405 132.470 ;
        RECT 163.405 130.195 175.405 130.220 ;
        RECT 176.730 132.470 177.680 135.495 ;
        RECT 187.805 135.470 188.730 135.495 ;
        RECT 178.455 132.470 179.255 135.470 ;
        RECT 179.755 132.470 180.555 135.470 ;
        RECT 176.730 132.445 177.655 132.470 ;
        RECT 176.730 130.220 177.480 132.445 ;
        RECT 177.730 132.080 178.690 132.310 ;
        RECT 178.830 132.195 179.255 132.470 ;
        RECT 181.030 132.195 181.830 135.470 ;
        RECT 182.330 132.470 183.130 135.470 ;
        RECT 183.605 132.195 184.405 135.470 ;
        RECT 184.905 132.470 185.705 135.470 ;
        RECT 186.180 132.470 186.980 135.470 ;
        RECT 187.770 132.470 188.730 135.470 ;
        RECT 186.180 132.195 186.605 132.470 ;
        RECT 177.730 130.670 178.580 132.080 ;
        RECT 178.830 131.395 186.605 132.195 ;
        RECT 186.760 132.080 187.720 132.310 ;
        RECT 178.930 130.220 186.505 131.020 ;
        RECT 186.855 130.670 187.705 132.080 ;
        RECT 187.955 130.220 188.730 132.470 ;
        RECT 176.730 130.195 188.730 130.220 ;
        RECT 190.055 132.445 191.005 135.470 ;
        RECT 191.780 132.470 192.580 135.470 ;
        RECT 193.080 132.470 193.880 135.470 ;
        RECT 190.055 130.195 190.780 132.445 ;
        RECT 191.055 132.080 192.015 132.310 ;
        RECT 192.155 132.195 192.580 132.470 ;
        RECT 194.355 132.195 195.155 135.470 ;
        RECT 195.630 132.470 196.430 135.470 ;
        RECT 196.930 132.470 197.730 135.470 ;
        RECT 198.515 132.470 199.480 135.470 ;
        RECT 196.930 132.195 197.355 132.470 ;
        RECT 198.530 132.445 199.480 132.470 ;
        RECT 191.055 130.670 191.905 132.080 ;
        RECT 192.155 131.395 197.355 132.195 ;
        RECT 197.505 132.080 198.465 132.310 ;
        RECT 192.255 130.195 197.255 131.120 ;
        RECT 197.555 130.670 198.405 132.080 ;
        RECT 198.680 130.195 199.480 132.445 ;
        RECT 200.805 132.470 201.755 135.495 ;
        RECT 211.880 135.470 212.805 135.495 ;
        RECT 202.530 132.470 203.330 135.470 ;
        RECT 203.830 132.470 204.630 135.470 ;
        RECT 200.805 132.445 201.730 132.470 ;
        RECT 200.805 130.220 201.555 132.445 ;
        RECT 201.805 132.080 202.765 132.310 ;
        RECT 202.905 132.195 203.330 132.470 ;
        RECT 205.105 132.195 205.905 135.470 ;
        RECT 206.405 132.470 207.205 135.470 ;
        RECT 207.680 132.195 208.480 135.470 ;
        RECT 208.980 132.470 209.780 135.470 ;
        RECT 210.255 132.470 211.055 135.470 ;
        RECT 211.845 132.470 212.805 135.470 ;
        RECT 210.255 132.195 210.680 132.470 ;
        RECT 201.805 130.670 202.655 132.080 ;
        RECT 202.905 131.395 210.680 132.195 ;
        RECT 210.835 132.080 211.795 132.310 ;
        RECT 203.005 130.220 210.580 131.020 ;
        RECT 210.930 130.670 211.780 132.080 ;
        RECT 212.030 130.220 212.805 132.470 ;
        RECT 200.805 130.195 212.805 130.220 ;
        RECT 214.130 132.470 215.080 135.495 ;
        RECT 225.205 135.470 228.050 135.495 ;
        RECT 215.855 132.470 216.655 135.470 ;
        RECT 217.155 132.470 217.955 135.470 ;
        RECT 214.130 132.445 215.055 132.470 ;
        RECT 214.130 130.220 214.880 132.445 ;
        RECT 215.130 132.080 216.090 132.310 ;
        RECT 216.230 132.195 216.655 132.470 ;
        RECT 218.430 132.195 219.230 135.470 ;
        RECT 219.730 132.470 220.530 135.470 ;
        RECT 221.005 132.195 221.805 135.470 ;
        RECT 222.305 132.470 223.105 135.470 ;
        RECT 223.580 132.470 224.380 135.470 ;
        RECT 225.170 132.470 228.050 135.470 ;
        RECT 223.580 132.195 224.005 132.470 ;
        RECT 215.130 130.670 215.980 132.080 ;
        RECT 216.230 131.395 224.005 132.195 ;
        RECT 224.160 132.080 225.120 132.310 ;
        RECT 216.330 130.220 223.905 131.020 ;
        RECT 224.255 130.670 225.105 132.080 ;
        RECT 225.355 130.220 228.050 132.470 ;
        RECT 214.130 130.195 228.050 130.220 ;
        RECT 75.025 129.450 228.050 130.195 ;
        RECT 75.030 129.445 228.050 129.450 ;
        RECT 111.950 128.135 113.050 128.250 ;
        RECT 97.830 128.100 98.080 128.135 ;
        RECT 98.660 128.100 98.910 128.135 ;
        RECT 99.490 128.100 99.740 128.135 ;
        RECT 100.320 128.100 100.570 128.135 ;
        RECT 101.150 128.100 101.400 128.135 ;
        RECT 101.980 128.100 102.230 128.135 ;
        RECT 102.810 128.100 103.060 128.135 ;
        RECT 103.640 128.100 103.890 128.135 ;
        RECT 104.470 128.100 104.720 128.135 ;
        RECT 105.300 128.100 105.550 128.135 ;
        RECT 106.130 128.100 106.380 128.135 ;
        RECT 106.960 128.100 107.210 128.135 ;
        RECT 107.790 128.100 108.040 128.135 ;
        RECT 108.620 128.100 108.870 128.135 ;
        RECT 109.450 128.100 109.700 128.135 ;
        RECT 110.280 128.100 110.530 128.135 ;
        RECT 111.110 128.100 111.360 128.135 ;
        RECT 47.925 126.075 98.100 128.100 ;
        RECT 98.650 126.075 99.750 128.100 ;
        RECT 100.320 126.075 101.425 128.100 ;
        RECT 101.975 126.075 103.075 128.100 ;
        RECT 103.640 126.075 104.750 128.100 ;
        RECT 105.300 126.075 106.400 128.100 ;
        RECT 106.960 126.075 108.075 128.100 ;
        RECT 108.620 126.075 109.725 128.100 ;
        RECT 110.275 126.075 111.375 128.100 ;
        RECT 111.940 127.200 113.050 128.135 ;
        RECT 111.925 126.075 113.050 127.200 ;
        RECT 113.600 128.100 113.850 128.135 ;
        RECT 114.430 128.100 114.680 128.135 ;
        RECT 115.260 128.100 115.510 128.135 ;
        RECT 116.090 128.100 116.340 128.135 ;
        RECT 116.920 128.100 117.170 128.135 ;
        RECT 117.750 128.100 118.000 128.135 ;
        RECT 118.580 128.100 118.830 128.135 ;
        RECT 119.410 128.100 119.660 128.135 ;
        RECT 120.240 128.100 120.490 128.135 ;
        RECT 121.070 128.100 121.320 128.135 ;
        RECT 121.900 128.100 122.150 128.135 ;
        RECT 122.730 128.100 122.980 128.135 ;
        RECT 123.560 128.100 123.810 128.135 ;
        RECT 124.390 128.100 124.640 128.135 ;
        RECT 125.220 128.100 125.470 128.135 ;
        RECT 126.050 128.100 126.300 128.135 ;
        RECT 126.880 128.100 127.130 128.135 ;
        RECT 127.710 128.100 127.960 128.135 ;
        RECT 128.540 128.100 128.790 128.135 ;
        RECT 129.370 128.100 129.620 128.135 ;
        RECT 130.200 128.100 130.450 128.135 ;
        RECT 131.030 128.100 131.280 128.135 ;
        RECT 131.860 128.100 132.110 128.135 ;
        RECT 132.690 128.100 132.940 128.135 ;
        RECT 133.520 128.100 133.770 128.135 ;
        RECT 134.350 128.100 134.600 128.135 ;
        RECT 135.180 128.100 135.430 128.135 ;
        RECT 136.010 128.100 136.260 128.135 ;
        RECT 136.840 128.100 137.090 128.135 ;
        RECT 137.670 128.100 137.920 128.135 ;
        RECT 138.500 128.100 138.750 128.135 ;
        RECT 139.330 128.100 139.580 128.135 ;
        RECT 140.160 128.100 140.410 128.135 ;
        RECT 140.990 128.100 141.240 128.135 ;
        RECT 141.820 128.100 142.070 128.135 ;
        RECT 142.650 128.100 142.900 128.135 ;
        RECT 143.480 128.100 143.730 128.135 ;
        RECT 144.310 128.100 144.560 128.135 ;
        RECT 145.140 128.100 145.390 128.135 ;
        RECT 145.970 128.100 146.220 128.135 ;
        RECT 146.800 128.100 147.050 128.135 ;
        RECT 147.630 128.100 147.880 128.135 ;
        RECT 148.460 128.100 148.710 128.135 ;
        RECT 149.290 128.100 149.540 128.135 ;
        RECT 150.120 128.100 150.370 128.135 ;
        RECT 150.950 128.100 151.200 128.135 ;
        RECT 151.780 128.100 152.030 128.135 ;
        RECT 152.610 128.100 152.860 128.135 ;
        RECT 153.440 128.100 153.690 128.135 ;
        RECT 154.270 128.100 154.520 128.135 ;
        RECT 155.100 128.100 155.350 128.135 ;
        RECT 155.930 128.100 156.180 128.135 ;
        RECT 156.760 128.100 157.010 128.135 ;
        RECT 157.590 128.100 157.840 128.135 ;
        RECT 158.420 128.100 158.670 128.135 ;
        RECT 159.250 128.100 159.500 128.135 ;
        RECT 160.080 128.100 160.330 128.135 ;
        RECT 160.910 128.100 161.160 128.135 ;
        RECT 161.740 128.100 161.990 128.135 ;
        RECT 162.570 128.100 162.820 128.135 ;
        RECT 163.400 128.100 163.650 128.135 ;
        RECT 164.230 128.100 164.480 128.135 ;
        RECT 165.060 128.100 165.310 128.135 ;
        RECT 165.890 128.100 166.140 128.135 ;
        RECT 166.720 128.100 166.970 128.135 ;
        RECT 167.550 128.100 167.800 128.135 ;
        RECT 168.380 128.100 168.630 128.135 ;
        RECT 169.210 128.100 169.460 128.135 ;
        RECT 170.040 128.100 170.290 128.135 ;
        RECT 170.870 128.100 171.120 128.135 ;
        RECT 171.700 128.100 171.950 128.135 ;
        RECT 172.530 128.100 172.780 128.135 ;
        RECT 173.360 128.100 173.610 128.135 ;
        RECT 174.190 128.100 174.440 128.135 ;
        RECT 175.020 128.100 175.270 128.135 ;
        RECT 175.850 128.100 176.100 128.135 ;
        RECT 176.680 128.100 176.930 128.135 ;
        RECT 177.510 128.100 177.760 128.135 ;
        RECT 178.340 128.100 178.590 128.135 ;
        RECT 179.170 128.100 179.420 128.135 ;
        RECT 113.600 126.075 114.700 128.100 ;
        RECT 115.260 126.075 116.375 128.100 ;
        RECT 116.920 126.075 118.025 128.100 ;
        RECT 118.575 126.075 119.675 128.100 ;
        RECT 120.240 126.075 121.350 128.100 ;
        RECT 121.900 126.075 123.000 128.100 ;
        RECT 123.560 126.075 124.675 128.100 ;
        RECT 125.220 126.075 126.325 128.100 ;
        RECT 126.880 126.075 128.000 128.100 ;
        RECT 128.540 126.075 129.650 128.100 ;
        RECT 130.200 126.075 131.300 128.100 ;
        RECT 131.860 126.075 132.975 128.100 ;
        RECT 133.520 126.075 134.625 128.100 ;
        RECT 135.175 126.075 136.275 128.100 ;
        RECT 136.840 126.075 137.950 128.100 ;
        RECT 138.500 126.075 139.600 128.100 ;
        RECT 140.160 126.075 141.275 128.100 ;
        RECT 141.820 126.075 142.925 128.100 ;
        RECT 143.475 126.075 144.575 128.100 ;
        RECT 145.125 126.075 146.225 128.100 ;
        RECT 146.800 126.075 147.900 128.100 ;
        RECT 148.460 126.075 149.575 128.100 ;
        RECT 150.120 126.075 151.225 128.100 ;
        RECT 151.775 126.075 152.875 128.100 ;
        RECT 153.440 126.075 154.550 128.100 ;
        RECT 155.100 126.075 156.200 128.100 ;
        RECT 156.750 126.075 157.850 128.100 ;
        RECT 158.420 126.075 159.525 128.100 ;
        RECT 160.075 126.075 161.175 128.100 ;
        RECT 161.740 126.075 162.850 128.100 ;
        RECT 163.400 126.075 164.500 128.100 ;
        RECT 165.060 126.075 166.175 128.100 ;
        RECT 166.720 126.075 167.825 128.100 ;
        RECT 168.375 126.075 169.475 128.100 ;
        RECT 170.040 126.075 171.150 128.100 ;
        RECT 171.700 126.075 172.800 128.100 ;
        RECT 173.360 126.075 174.475 128.100 ;
        RECT 175.020 126.075 176.125 128.100 ;
        RECT 176.675 126.075 177.775 128.100 ;
        RECT 178.340 126.075 179.450 128.100 ;
        RECT 47.925 12.775 49.950 126.075 ;
        RECT 97.830 126.030 98.080 126.075 ;
        RECT 98.660 126.030 98.910 126.075 ;
        RECT 99.490 126.030 99.740 126.075 ;
        RECT 100.320 126.030 100.570 126.075 ;
        RECT 101.150 126.030 101.400 126.075 ;
        RECT 101.980 126.030 102.230 126.075 ;
        RECT 102.810 126.030 103.060 126.075 ;
        RECT 103.640 126.030 103.890 126.075 ;
        RECT 104.470 126.030 104.720 126.075 ;
        RECT 105.300 126.030 105.550 126.075 ;
        RECT 106.130 126.030 106.380 126.075 ;
        RECT 106.960 126.030 107.210 126.075 ;
        RECT 107.790 126.030 108.040 126.075 ;
        RECT 108.620 126.030 108.870 126.075 ;
        RECT 109.450 126.030 109.700 126.075 ;
        RECT 110.280 126.030 110.530 126.075 ;
        RECT 111.110 126.030 111.360 126.075 ;
        RECT 111.940 126.030 112.190 126.075 ;
        RECT 112.770 126.030 113.020 126.075 ;
        RECT 113.600 126.030 113.850 126.075 ;
        RECT 114.430 126.030 114.680 126.075 ;
        RECT 115.260 126.030 115.510 126.075 ;
        RECT 116.090 126.030 116.340 126.075 ;
        RECT 116.920 126.030 117.170 126.075 ;
        RECT 117.750 126.030 118.000 126.075 ;
        RECT 118.580 126.030 118.830 126.075 ;
        RECT 119.410 126.030 119.660 126.075 ;
        RECT 120.240 126.030 120.490 126.075 ;
        RECT 121.070 126.030 121.320 126.075 ;
        RECT 121.900 126.030 122.150 126.075 ;
        RECT 122.730 126.030 122.980 126.075 ;
        RECT 123.560 126.030 123.810 126.075 ;
        RECT 124.390 126.030 124.640 126.075 ;
        RECT 125.220 126.030 125.470 126.075 ;
        RECT 126.050 126.030 126.300 126.075 ;
        RECT 126.880 126.030 127.130 126.075 ;
        RECT 127.710 126.030 127.960 126.075 ;
        RECT 128.540 126.030 128.790 126.075 ;
        RECT 129.370 126.030 129.620 126.075 ;
        RECT 130.200 126.030 130.450 126.075 ;
        RECT 131.030 126.030 131.280 126.075 ;
        RECT 131.860 126.030 132.110 126.075 ;
        RECT 132.690 126.030 132.940 126.075 ;
        RECT 133.520 126.030 133.770 126.075 ;
        RECT 134.350 126.030 134.600 126.075 ;
        RECT 135.180 126.030 135.430 126.075 ;
        RECT 136.010 126.030 136.260 126.075 ;
        RECT 136.840 126.030 137.090 126.075 ;
        RECT 137.670 126.030 137.920 126.075 ;
        RECT 138.500 126.030 138.750 126.075 ;
        RECT 139.330 126.030 139.580 126.075 ;
        RECT 140.160 126.030 140.410 126.075 ;
        RECT 140.990 126.030 141.240 126.075 ;
        RECT 141.820 126.030 142.070 126.075 ;
        RECT 142.650 126.030 142.900 126.075 ;
        RECT 143.480 126.030 143.730 126.075 ;
        RECT 144.310 126.030 144.560 126.075 ;
        RECT 145.140 126.030 145.390 126.075 ;
        RECT 145.970 126.030 146.220 126.075 ;
        RECT 146.800 126.030 147.050 126.075 ;
        RECT 147.630 126.030 147.880 126.075 ;
        RECT 148.460 126.030 148.710 126.075 ;
        RECT 149.290 126.030 149.540 126.075 ;
        RECT 150.120 126.030 150.370 126.075 ;
        RECT 150.950 126.030 151.200 126.075 ;
        RECT 151.780 126.030 152.030 126.075 ;
        RECT 152.610 126.030 152.860 126.075 ;
        RECT 153.440 126.030 153.690 126.075 ;
        RECT 154.270 126.030 154.520 126.075 ;
        RECT 155.100 126.030 155.350 126.075 ;
        RECT 155.930 126.030 156.180 126.075 ;
        RECT 156.760 126.030 157.010 126.075 ;
        RECT 157.590 126.030 157.840 126.075 ;
        RECT 158.420 126.030 158.670 126.075 ;
        RECT 159.250 126.030 159.500 126.075 ;
        RECT 160.080 126.030 160.330 126.075 ;
        RECT 160.910 126.030 161.160 126.075 ;
        RECT 161.740 126.030 161.990 126.075 ;
        RECT 162.570 126.030 162.820 126.075 ;
        RECT 163.400 126.030 163.650 126.075 ;
        RECT 164.230 126.030 164.480 126.075 ;
        RECT 165.060 126.030 165.310 126.075 ;
        RECT 165.890 126.030 166.140 126.075 ;
        RECT 166.720 126.030 166.970 126.075 ;
        RECT 167.550 126.030 167.800 126.075 ;
        RECT 168.380 126.030 168.630 126.075 ;
        RECT 169.210 126.030 169.460 126.075 ;
        RECT 170.040 126.030 170.290 126.075 ;
        RECT 170.870 126.030 171.120 126.075 ;
        RECT 171.700 126.030 171.950 126.075 ;
        RECT 172.530 126.030 172.780 126.075 ;
        RECT 173.360 126.030 173.610 126.075 ;
        RECT 174.190 126.030 174.440 126.075 ;
        RECT 175.020 126.030 175.270 126.075 ;
        RECT 175.850 126.030 176.100 126.075 ;
        RECT 176.680 126.030 176.930 126.075 ;
        RECT 177.510 126.030 177.760 126.075 ;
        RECT 178.340 126.030 178.590 126.075 ;
        RECT 179.170 126.030 179.420 126.075 ;
        RECT 179.900 126.025 180.350 128.150 ;
        RECT 180.650 126.025 181.250 128.150 ;
        RECT 181.660 128.100 181.910 128.135 ;
        RECT 182.490 128.100 182.740 128.135 ;
        RECT 183.320 128.100 183.570 128.135 ;
        RECT 184.150 128.100 184.400 128.135 ;
        RECT 184.980 128.100 185.230 128.135 ;
        RECT 185.810 128.100 186.060 128.135 ;
        RECT 186.640 128.100 186.890 128.135 ;
        RECT 187.470 128.100 187.720 128.135 ;
        RECT 188.300 128.100 188.550 128.135 ;
        RECT 189.130 128.100 189.380 128.135 ;
        RECT 189.960 128.100 190.210 128.135 ;
        RECT 190.790 128.100 191.040 128.135 ;
        RECT 191.620 128.100 191.870 128.135 ;
        RECT 192.450 128.100 192.700 128.135 ;
        RECT 193.280 128.100 193.530 128.135 ;
        RECT 194.110 128.100 194.360 128.135 ;
        RECT 194.940 128.100 195.190 128.135 ;
        RECT 195.770 128.100 196.020 128.135 ;
        RECT 196.600 128.100 196.850 128.135 ;
        RECT 197.430 128.100 197.680 128.135 ;
        RECT 198.260 128.100 198.510 128.135 ;
        RECT 199.090 128.100 199.340 128.135 ;
        RECT 199.920 128.100 200.170 128.135 ;
        RECT 200.750 128.100 201.000 128.135 ;
        RECT 201.580 128.100 201.830 128.135 ;
        RECT 202.410 128.100 202.660 128.135 ;
        RECT 203.240 128.100 203.490 128.135 ;
        RECT 204.070 128.100 204.320 128.135 ;
        RECT 204.900 128.100 205.150 128.135 ;
        RECT 205.730 128.100 205.980 128.135 ;
        RECT 206.560 128.100 206.810 128.135 ;
        RECT 207.390 128.100 207.640 128.135 ;
        RECT 208.220 128.100 208.470 128.135 ;
        RECT 209.050 128.100 209.300 128.135 ;
        RECT 209.880 128.100 210.130 128.135 ;
        RECT 210.710 128.100 210.960 128.135 ;
        RECT 211.540 128.100 211.790 128.135 ;
        RECT 181.660 126.075 182.775 128.100 ;
        RECT 183.320 126.075 184.425 128.100 ;
        RECT 184.975 126.075 186.075 128.100 ;
        RECT 186.640 126.075 187.750 128.100 ;
        RECT 188.300 126.075 189.400 128.100 ;
        RECT 189.960 126.075 191.075 128.100 ;
        RECT 191.620 126.075 192.725 128.100 ;
        RECT 193.275 126.075 194.375 128.100 ;
        RECT 194.940 126.075 196.050 128.100 ;
        RECT 196.600 126.075 197.700 128.100 ;
        RECT 198.260 126.075 199.375 128.100 ;
        RECT 199.920 126.075 201.025 128.100 ;
        RECT 201.575 126.075 202.675 128.100 ;
        RECT 203.240 126.075 204.350 128.100 ;
        RECT 204.900 126.075 206.000 128.100 ;
        RECT 206.560 126.075 207.675 128.100 ;
        RECT 208.220 126.075 209.325 128.100 ;
        RECT 209.875 126.075 210.975 128.100 ;
        RECT 211.540 126.075 214.125 128.100 ;
        RECT 181.660 126.030 181.910 126.075 ;
        RECT 182.490 126.030 182.740 126.075 ;
        RECT 183.320 126.030 183.570 126.075 ;
        RECT 184.150 126.030 184.400 126.075 ;
        RECT 184.980 126.030 185.230 126.075 ;
        RECT 185.810 126.030 186.060 126.075 ;
        RECT 186.640 126.030 186.890 126.075 ;
        RECT 187.470 126.030 187.720 126.075 ;
        RECT 188.300 126.030 188.550 126.075 ;
        RECT 189.130 126.030 189.380 126.075 ;
        RECT 189.960 126.030 190.210 126.075 ;
        RECT 190.790 126.030 191.040 126.075 ;
        RECT 191.620 126.030 191.870 126.075 ;
        RECT 192.450 126.030 192.700 126.075 ;
        RECT 193.280 126.030 193.530 126.075 ;
        RECT 194.110 126.030 194.360 126.075 ;
        RECT 194.940 126.030 195.190 126.075 ;
        RECT 195.770 126.030 196.020 126.075 ;
        RECT 196.600 126.030 196.850 126.075 ;
        RECT 197.430 126.030 197.680 126.075 ;
        RECT 198.260 126.030 198.510 126.075 ;
        RECT 199.090 126.030 199.340 126.075 ;
        RECT 199.920 126.030 200.170 126.075 ;
        RECT 200.750 126.030 201.000 126.075 ;
        RECT 201.580 126.030 201.830 126.075 ;
        RECT 202.410 126.030 202.660 126.075 ;
        RECT 203.240 126.030 203.490 126.075 ;
        RECT 204.070 126.030 204.320 126.075 ;
        RECT 204.900 126.030 205.150 126.075 ;
        RECT 205.730 126.030 205.980 126.075 ;
        RECT 206.560 126.030 206.810 126.075 ;
        RECT 207.390 126.030 207.640 126.075 ;
        RECT 208.220 126.030 208.470 126.075 ;
        RECT 209.050 126.030 209.300 126.075 ;
        RECT 209.880 126.030 210.130 126.075 ;
        RECT 210.710 126.030 210.960 126.075 ;
        RECT 211.540 126.030 211.790 126.075 ;
        RECT 215.625 125.400 228.050 129.445 ;
        RECT 75.275 121.525 97.300 125.400 ;
        RECT 97.830 124.100 98.080 124.140 ;
        RECT 98.660 124.100 98.910 124.140 ;
        RECT 99.490 124.100 99.740 124.140 ;
        RECT 100.320 124.100 100.570 124.140 ;
        RECT 101.150 124.100 101.400 124.140 ;
        RECT 101.980 124.100 102.230 124.140 ;
        RECT 102.810 124.100 103.060 124.140 ;
        RECT 103.640 124.100 103.890 124.140 ;
        RECT 104.470 124.100 104.720 124.140 ;
        RECT 105.300 124.100 105.550 124.140 ;
        RECT 106.130 124.100 106.380 124.140 ;
        RECT 106.960 124.100 107.210 124.140 ;
        RECT 107.790 124.100 108.040 124.140 ;
        RECT 108.620 124.100 108.870 124.140 ;
        RECT 109.450 124.100 109.700 124.140 ;
        RECT 110.280 124.100 110.530 124.140 ;
        RECT 111.110 124.100 111.360 124.140 ;
        RECT 111.940 124.100 112.190 124.140 ;
        RECT 112.770 124.100 113.020 124.140 ;
        RECT 113.600 124.100 113.850 124.140 ;
        RECT 114.430 124.100 114.680 124.140 ;
        RECT 115.260 124.100 115.510 124.140 ;
        RECT 116.090 124.100 116.340 124.140 ;
        RECT 116.920 124.100 117.170 124.140 ;
        RECT 117.750 124.100 118.000 124.140 ;
        RECT 118.580 124.100 118.830 124.140 ;
        RECT 119.410 124.100 119.660 124.140 ;
        RECT 120.240 124.100 120.490 124.140 ;
        RECT 121.070 124.100 121.320 124.140 ;
        RECT 121.900 124.100 122.150 124.140 ;
        RECT 122.730 124.100 122.980 124.140 ;
        RECT 123.560 124.100 123.810 124.140 ;
        RECT 124.390 124.100 124.640 124.140 ;
        RECT 125.220 124.100 125.470 124.140 ;
        RECT 126.050 124.100 126.300 124.140 ;
        RECT 126.880 124.100 127.130 124.140 ;
        RECT 97.825 122.075 98.925 124.100 ;
        RECT 99.475 122.075 100.600 124.100 ;
        RECT 101.150 122.075 102.250 124.100 ;
        RECT 102.800 122.075 103.900 124.100 ;
        RECT 104.470 122.075 105.575 124.100 ;
        RECT 106.125 122.075 107.225 124.100 ;
        RECT 107.775 122.075 108.875 124.100 ;
        RECT 109.450 122.075 110.550 124.100 ;
        RECT 111.100 122.075 112.200 124.100 ;
        RECT 112.770 122.075 113.875 124.100 ;
        RECT 114.425 122.075 115.525 124.100 ;
        RECT 116.090 122.075 117.200 124.100 ;
        RECT 117.750 122.075 118.850 124.100 ;
        RECT 119.400 122.075 120.500 124.100 ;
        RECT 121.070 122.075 122.175 124.100 ;
        RECT 122.725 122.075 123.825 124.100 ;
        RECT 124.390 122.075 125.500 124.100 ;
        RECT 126.050 122.075 127.150 124.100 ;
        RECT 97.830 122.035 98.080 122.075 ;
        RECT 98.660 122.035 98.910 122.075 ;
        RECT 99.490 122.035 99.740 122.075 ;
        RECT 100.320 122.035 100.570 122.075 ;
        RECT 101.150 122.035 101.400 122.075 ;
        RECT 101.980 122.035 102.230 122.075 ;
        RECT 102.810 122.035 103.060 122.075 ;
        RECT 103.640 122.035 103.890 122.075 ;
        RECT 104.470 122.035 104.720 122.075 ;
        RECT 105.300 122.035 105.550 122.075 ;
        RECT 106.130 122.035 106.380 122.075 ;
        RECT 106.960 122.035 107.210 122.075 ;
        RECT 107.790 122.035 108.040 122.075 ;
        RECT 108.620 122.035 108.870 122.075 ;
        RECT 109.450 122.035 109.700 122.075 ;
        RECT 110.280 122.035 110.530 122.075 ;
        RECT 111.110 122.035 111.360 122.075 ;
        RECT 111.940 122.035 112.190 122.075 ;
        RECT 112.770 122.035 113.020 122.075 ;
        RECT 113.600 122.035 113.850 122.075 ;
        RECT 114.430 122.035 114.680 122.075 ;
        RECT 115.260 122.035 115.510 122.075 ;
        RECT 116.090 122.035 116.340 122.075 ;
        RECT 116.920 122.035 117.170 122.075 ;
        RECT 117.750 122.035 118.000 122.075 ;
        RECT 118.580 122.035 118.830 122.075 ;
        RECT 119.410 122.035 119.660 122.075 ;
        RECT 120.240 122.035 120.490 122.075 ;
        RECT 121.070 122.035 121.320 122.075 ;
        RECT 121.900 122.035 122.150 122.075 ;
        RECT 122.730 122.035 122.980 122.075 ;
        RECT 123.560 122.035 123.810 122.075 ;
        RECT 124.390 122.035 124.640 122.075 ;
        RECT 125.220 122.035 125.470 122.075 ;
        RECT 126.050 122.035 126.300 122.075 ;
        RECT 126.880 122.035 127.130 122.075 ;
        RECT 127.675 122.025 128.825 124.150 ;
        RECT 129.370 124.100 129.620 124.140 ;
        RECT 130.200 124.100 130.450 124.140 ;
        RECT 131.030 124.100 131.280 124.140 ;
        RECT 131.860 124.100 132.110 124.140 ;
        RECT 132.690 124.100 132.940 124.140 ;
        RECT 133.520 124.100 133.770 124.140 ;
        RECT 134.350 124.100 134.600 124.140 ;
        RECT 135.180 124.100 135.430 124.140 ;
        RECT 136.010 124.100 136.260 124.140 ;
        RECT 136.840 124.100 137.090 124.140 ;
        RECT 137.670 124.100 137.920 124.140 ;
        RECT 138.500 124.100 138.750 124.140 ;
        RECT 139.330 124.100 139.580 124.140 ;
        RECT 140.160 124.100 140.410 124.140 ;
        RECT 140.990 124.100 141.240 124.140 ;
        RECT 141.820 124.100 142.070 124.140 ;
        RECT 142.650 124.100 142.900 124.140 ;
        RECT 143.480 124.100 143.730 124.140 ;
        RECT 144.310 124.100 144.560 124.140 ;
        RECT 145.140 124.100 145.390 124.140 ;
        RECT 145.970 124.100 146.220 124.140 ;
        RECT 146.800 124.100 147.050 124.140 ;
        RECT 147.630 124.100 147.880 124.140 ;
        RECT 148.460 124.100 148.710 124.140 ;
        RECT 149.290 124.100 149.540 124.140 ;
        RECT 150.120 124.100 150.370 124.140 ;
        RECT 150.950 124.100 151.200 124.140 ;
        RECT 151.780 124.100 152.030 124.140 ;
        RECT 152.610 124.100 152.860 124.140 ;
        RECT 153.440 124.100 153.690 124.140 ;
        RECT 154.270 124.100 154.520 124.140 ;
        RECT 155.100 124.100 155.350 124.140 ;
        RECT 155.930 124.100 156.180 124.140 ;
        RECT 156.760 124.100 157.010 124.140 ;
        RECT 157.590 124.100 157.840 124.140 ;
        RECT 158.420 124.100 158.670 124.140 ;
        RECT 159.250 124.100 159.500 124.140 ;
        RECT 160.080 124.100 160.330 124.140 ;
        RECT 160.910 124.100 161.160 124.140 ;
        RECT 161.740 124.100 161.990 124.140 ;
        RECT 162.570 124.100 162.820 124.140 ;
        RECT 163.400 124.100 163.650 124.140 ;
        RECT 164.230 124.100 164.480 124.140 ;
        RECT 165.060 124.100 165.310 124.140 ;
        RECT 165.890 124.100 166.140 124.140 ;
        RECT 166.720 124.100 166.970 124.140 ;
        RECT 167.550 124.100 167.800 124.140 ;
        RECT 168.380 124.100 168.630 124.140 ;
        RECT 169.210 124.100 169.460 124.140 ;
        RECT 170.040 124.100 170.290 124.140 ;
        RECT 170.870 124.100 171.120 124.140 ;
        RECT 171.700 124.100 171.950 124.140 ;
        RECT 172.530 124.100 172.780 124.140 ;
        RECT 173.360 124.100 173.610 124.140 ;
        RECT 174.190 124.100 174.440 124.140 ;
        RECT 175.020 124.100 175.270 124.140 ;
        RECT 175.850 124.100 176.100 124.140 ;
        RECT 176.680 124.100 176.930 124.140 ;
        RECT 177.510 124.100 177.760 124.140 ;
        RECT 178.340 124.100 178.590 124.140 ;
        RECT 179.170 124.100 179.420 124.140 ;
        RECT 180.000 124.100 180.250 124.140 ;
        RECT 180.830 124.100 181.080 124.140 ;
        RECT 181.660 124.100 181.910 124.140 ;
        RECT 182.490 124.100 182.740 124.140 ;
        RECT 183.320 124.100 183.570 124.140 ;
        RECT 184.150 124.100 184.400 124.140 ;
        RECT 184.980 124.100 185.230 124.140 ;
        RECT 185.810 124.100 186.060 124.140 ;
        RECT 186.640 124.100 186.890 124.140 ;
        RECT 187.470 124.100 187.720 124.140 ;
        RECT 188.300 124.100 188.550 124.140 ;
        RECT 189.130 124.100 189.380 124.140 ;
        RECT 189.960 124.100 190.210 124.140 ;
        RECT 190.790 124.100 191.040 124.140 ;
        RECT 191.620 124.100 191.870 124.140 ;
        RECT 192.450 124.100 192.700 124.140 ;
        RECT 193.280 124.100 193.530 124.140 ;
        RECT 194.110 124.100 194.360 124.140 ;
        RECT 194.940 124.100 195.190 124.140 ;
        RECT 195.770 124.100 196.020 124.140 ;
        RECT 196.600 124.100 196.850 124.140 ;
        RECT 197.430 124.100 197.680 124.140 ;
        RECT 198.260 124.100 198.510 124.140 ;
        RECT 199.090 124.100 199.340 124.140 ;
        RECT 199.920 124.100 200.170 124.140 ;
        RECT 200.750 124.100 201.000 124.140 ;
        RECT 201.580 124.100 201.830 124.140 ;
        RECT 202.410 124.100 202.660 124.140 ;
        RECT 203.240 124.100 203.490 124.140 ;
        RECT 204.070 124.100 204.320 124.140 ;
        RECT 204.900 124.100 205.150 124.140 ;
        RECT 205.730 124.100 205.980 124.140 ;
        RECT 206.560 124.100 206.810 124.140 ;
        RECT 207.390 124.100 207.640 124.140 ;
        RECT 208.220 124.100 208.470 124.140 ;
        RECT 209.050 124.100 209.300 124.140 ;
        RECT 209.880 124.100 210.130 124.140 ;
        RECT 210.710 124.100 210.960 124.140 ;
        RECT 211.540 124.100 211.790 124.140 ;
        RECT 129.370 122.075 130.475 124.100 ;
        RECT 131.025 122.075 132.125 124.100 ;
        RECT 132.690 122.075 133.800 124.100 ;
        RECT 134.350 122.075 135.450 124.100 ;
        RECT 136.000 122.075 137.100 124.100 ;
        RECT 137.670 122.075 138.775 124.100 ;
        RECT 139.325 122.075 140.425 124.100 ;
        RECT 140.990 122.075 142.100 124.100 ;
        RECT 142.650 122.075 143.750 124.100 ;
        RECT 144.310 122.075 145.425 124.100 ;
        RECT 145.970 122.075 147.075 124.100 ;
        RECT 147.625 122.075 148.725 124.100 ;
        RECT 149.290 122.075 150.400 124.100 ;
        RECT 150.950 122.075 152.050 124.100 ;
        RECT 152.610 122.075 153.725 124.100 ;
        RECT 154.270 122.075 155.375 124.100 ;
        RECT 155.925 122.075 157.025 124.100 ;
        RECT 157.590 122.075 158.700 124.100 ;
        RECT 159.250 122.075 160.350 124.100 ;
        RECT 160.900 122.075 162.000 124.100 ;
        RECT 162.570 122.075 163.675 124.100 ;
        RECT 164.225 122.075 165.325 124.100 ;
        RECT 165.890 122.075 167.000 124.100 ;
        RECT 167.550 122.075 168.650 124.100 ;
        RECT 169.200 122.075 170.300 124.100 ;
        RECT 170.850 122.075 171.950 124.100 ;
        RECT 172.525 122.075 173.625 124.100 ;
        RECT 174.190 122.075 175.300 124.100 ;
        RECT 175.850 122.075 176.950 124.100 ;
        RECT 177.500 122.075 178.600 124.100 ;
        RECT 179.170 122.075 180.275 124.100 ;
        RECT 180.825 122.075 181.925 124.100 ;
        RECT 182.490 122.075 183.600 124.100 ;
        RECT 184.150 122.075 185.250 124.100 ;
        RECT 185.810 122.075 186.925 124.100 ;
        RECT 187.470 122.075 188.575 124.100 ;
        RECT 189.125 122.075 190.225 124.100 ;
        RECT 190.775 122.075 191.875 124.100 ;
        RECT 192.450 122.075 193.550 124.100 ;
        RECT 194.100 122.075 195.200 124.100 ;
        RECT 195.750 122.075 196.850 124.100 ;
        RECT 197.425 122.075 198.525 124.100 ;
        RECT 199.090 122.075 200.200 124.100 ;
        RECT 200.750 122.075 201.850 124.100 ;
        RECT 202.400 122.075 203.500 124.100 ;
        RECT 204.070 122.075 205.175 124.100 ;
        RECT 205.725 122.075 206.825 124.100 ;
        RECT 207.375 122.075 208.475 124.100 ;
        RECT 209.050 122.075 210.150 124.100 ;
        RECT 210.700 122.075 211.800 124.100 ;
        RECT 212.325 122.350 228.050 125.400 ;
        RECT 230.000 133.125 230.600 139.800 ;
        RECT 231.050 138.145 266.400 139.000 ;
        RECT 231.045 137.800 266.400 138.145 ;
        RECT 231.045 137.795 234.650 137.800 ;
        RECT 235.645 137.795 248.450 137.800 ;
        RECT 231.050 137.775 234.650 137.795 ;
        RECT 231.050 137.050 232.050 137.775 ;
        RECT 233.650 137.595 234.650 137.775 ;
        RECT 233.645 137.270 234.650 137.595 ;
        RECT 233.650 137.050 234.650 137.270 ;
        RECT 231.050 137.045 232.275 137.050 ;
        RECT 231.050 134.050 232.480 137.045 ;
        RECT 232.675 134.050 233.025 137.050 ;
        RECT 233.425 137.045 234.650 137.050 ;
        RECT 233.210 134.050 234.650 137.045 ;
        RECT 235.650 137.775 248.450 137.795 ;
        RECT 235.650 137.050 236.650 137.775 ;
        RECT 238.250 137.595 241.525 137.775 ;
        RECT 242.575 137.595 245.850 137.775 ;
        RECT 247.450 137.595 248.450 137.775 ;
        RECT 238.245 137.275 241.525 137.595 ;
        RECT 238.245 137.270 241.250 137.275 ;
        RECT 242.570 137.270 245.850 137.595 ;
        RECT 247.445 137.270 248.450 137.595 ;
        RECT 238.250 137.050 241.250 137.270 ;
        RECT 242.850 137.050 245.850 137.270 ;
        RECT 247.450 137.050 248.450 137.270 ;
        RECT 235.650 137.045 236.875 137.050 ;
        RECT 235.650 134.050 237.080 137.045 ;
        RECT 237.275 134.050 237.625 137.050 ;
        RECT 238.025 137.045 241.475 137.050 ;
        RECT 237.810 134.050 241.680 137.045 ;
        RECT 241.875 134.050 242.225 137.050 ;
        RECT 242.625 137.045 246.075 137.050 ;
        RECT 242.410 134.050 246.280 137.045 ;
        RECT 246.475 134.050 246.825 137.050 ;
        RECT 247.225 137.045 248.450 137.050 ;
        RECT 247.010 134.050 248.450 137.045 ;
        RECT 249.450 137.600 250.450 137.800 ;
        RECT 249.450 137.275 250.455 137.600 ;
        RECT 249.450 137.050 250.450 137.275 ;
        RECT 249.450 134.050 250.880 137.050 ;
        RECT 251.075 134.050 251.400 137.050 ;
        RECT 251.600 134.050 251.850 137.800 ;
        RECT 252.050 134.050 252.375 137.050 ;
        RECT 252.550 134.050 252.800 137.800 ;
        RECT 253.950 137.650 266.400 137.800 ;
        RECT 253.950 137.050 254.950 137.650 ;
        RECT 253.000 134.050 253.325 137.050 ;
        RECT 253.530 134.050 254.950 137.050 ;
        RECT 231.770 134.045 232.000 134.050 ;
        RECT 232.250 134.045 232.480 134.050 ;
        RECT 232.730 134.045 232.960 134.050 ;
        RECT 233.210 134.045 233.440 134.050 ;
        RECT 233.690 134.045 233.920 134.050 ;
        RECT 236.370 134.045 236.600 134.050 ;
        RECT 236.850 134.045 237.080 134.050 ;
        RECT 237.330 134.045 237.560 134.050 ;
        RECT 237.810 134.045 238.040 134.050 ;
        RECT 238.290 134.045 238.520 134.050 ;
        RECT 240.970 134.045 241.200 134.050 ;
        RECT 241.450 134.045 241.680 134.050 ;
        RECT 241.930 134.045 242.160 134.050 ;
        RECT 242.410 134.045 242.640 134.050 ;
        RECT 242.890 134.045 243.120 134.050 ;
        RECT 245.570 134.045 245.800 134.050 ;
        RECT 246.050 134.045 246.280 134.050 ;
        RECT 246.530 134.045 246.760 134.050 ;
        RECT 247.010 134.045 247.240 134.050 ;
        RECT 247.490 134.045 247.720 134.050 ;
        RECT 232.450 133.845 233.250 133.850 ;
        RECT 237.050 133.845 237.850 133.850 ;
        RECT 242.100 133.845 242.475 133.850 ;
        RECT 246.250 133.845 247.050 133.850 ;
        RECT 232.445 133.470 233.250 133.845 ;
        RECT 237.045 133.470 237.850 133.845 ;
        RECT 242.095 133.470 242.475 133.845 ;
        RECT 246.245 133.470 247.050 133.845 ;
        RECT 232.450 133.125 233.250 133.470 ;
        RECT 237.050 133.125 237.850 133.470 ;
        RECT 242.100 133.125 242.475 133.470 ;
        RECT 246.250 133.125 247.050 133.470 ;
        RECT 250.825 133.475 253.580 133.850 ;
        RECT 250.825 133.125 253.575 133.475 ;
        RECT 230.000 132.525 233.250 133.125 ;
        RECT 234.900 132.525 237.850 133.125 ;
        RECT 239.500 132.525 242.475 133.125 ;
        RECT 244.775 132.525 247.050 133.125 ;
        RECT 248.700 132.525 253.575 133.125 ;
        RECT 230.000 123.825 230.600 132.525 ;
        RECT 232.450 131.850 233.250 132.525 ;
        RECT 237.050 131.850 237.850 132.525 ;
        RECT 242.100 131.850 242.475 132.525 ;
        RECT 246.250 131.850 247.050 132.525 ;
        RECT 250.825 132.175 253.575 132.525 ;
        RECT 250.825 131.850 253.580 132.175 ;
        RECT 256.625 132.100 271.250 132.450 ;
        RECT 231.050 130.650 232.485 131.650 ;
        RECT 232.675 130.650 233.025 131.650 ;
        RECT 233.215 130.650 237.085 131.650 ;
        RECT 237.275 130.650 237.625 131.650 ;
        RECT 237.815 130.650 239.250 131.650 ;
        RECT 231.050 129.950 232.050 130.650 ;
        RECT 233.650 129.950 236.650 130.650 ;
        RECT 238.250 129.950 239.250 130.650 ;
        RECT 240.250 130.650 241.685 131.650 ;
        RECT 241.875 130.650 242.225 131.650 ;
        RECT 242.415 130.650 243.850 131.650 ;
        RECT 240.250 130.450 241.250 130.650 ;
        RECT 242.850 130.450 243.850 130.650 ;
        RECT 240.250 129.950 241.525 130.450 ;
        RECT 242.575 129.950 243.850 130.450 ;
        RECT 244.850 130.650 246.285 131.650 ;
        RECT 246.475 130.650 246.825 131.650 ;
        RECT 247.015 130.650 250.880 131.650 ;
        RECT 251.075 130.650 251.400 131.650 ;
        RECT 244.850 129.950 245.850 130.650 ;
        RECT 247.450 130.625 250.880 130.650 ;
        RECT 247.450 129.950 250.875 130.625 ;
        RECT 251.600 129.950 251.850 131.650 ;
        RECT 252.050 130.650 252.375 131.650 ;
        RECT 252.550 129.950 252.800 131.650 ;
        RECT 253.000 130.650 253.325 131.650 ;
        RECT 253.525 129.950 254.950 131.650 ;
        RECT 256.625 131.550 271.250 131.925 ;
        RECT 231.050 129.600 254.955 129.950 ;
        RECT 231.050 128.850 233.700 128.855 ;
        RECT 231.050 128.500 254.955 128.850 ;
        RECT 231.050 124.750 231.425 128.500 ;
        RECT 231.950 127.950 232.800 128.330 ;
        RECT 231.775 123.825 232.025 127.775 ;
        RECT 232.200 124.750 232.550 127.775 ;
        RECT 232.725 123.825 232.975 127.775 ;
        RECT 233.325 124.750 233.700 128.500 ;
        RECT 235.645 128.495 248.450 128.500 ;
        RECT 235.650 128.475 248.450 128.495 ;
        RECT 235.650 127.750 236.650 128.475 ;
        RECT 238.250 128.295 241.525 128.475 ;
        RECT 242.575 128.295 245.850 128.475 ;
        RECT 247.450 128.295 248.450 128.475 ;
        RECT 238.245 127.975 241.525 128.295 ;
        RECT 238.245 127.970 241.250 127.975 ;
        RECT 242.570 127.970 245.850 128.295 ;
        RECT 247.445 127.970 248.450 128.295 ;
        RECT 238.250 127.750 241.250 127.970 ;
        RECT 242.850 127.750 245.850 127.970 ;
        RECT 247.450 127.750 248.450 127.970 ;
        RECT 235.650 127.745 236.875 127.750 ;
        RECT 235.650 124.750 237.080 127.745 ;
        RECT 237.275 124.750 237.625 127.750 ;
        RECT 238.025 127.745 241.475 127.750 ;
        RECT 237.810 124.750 241.680 127.745 ;
        RECT 241.875 124.750 242.225 127.750 ;
        RECT 242.625 127.745 246.075 127.750 ;
        RECT 242.410 124.750 246.280 127.745 ;
        RECT 246.475 124.750 246.825 127.750 ;
        RECT 247.225 127.745 248.450 127.750 ;
        RECT 247.010 124.750 248.450 127.745 ;
        RECT 249.450 128.300 250.450 128.500 ;
        RECT 249.450 127.975 250.455 128.300 ;
        RECT 249.450 127.750 250.450 127.975 ;
        RECT 249.450 124.750 250.880 127.750 ;
        RECT 251.075 124.750 251.400 127.750 ;
        RECT 251.600 124.750 251.850 128.500 ;
        RECT 252.050 124.750 252.375 127.750 ;
        RECT 252.550 124.750 252.800 128.500 ;
        RECT 253.950 127.750 254.950 128.500 ;
        RECT 253.000 124.750 253.325 127.750 ;
        RECT 253.530 124.750 254.950 127.750 ;
        RECT 256.625 124.750 256.975 131.550 ;
        RECT 257.540 131.545 259.290 131.550 ;
        RECT 268.590 131.545 270.340 131.550 ;
        RECT 257.345 131.275 257.575 131.345 ;
        RECT 257.825 131.275 258.055 131.345 ;
        RECT 258.305 131.275 258.535 131.345 ;
        RECT 258.785 131.275 259.015 131.345 ;
        RECT 259.265 131.275 259.495 131.345 ;
        RECT 259.745 131.275 259.975 131.345 ;
        RECT 257.300 130.100 259.500 131.275 ;
        RECT 259.700 130.100 260.025 131.275 ;
        RECT 257.345 128.345 257.575 130.100 ;
        RECT 257.825 128.345 258.055 130.100 ;
        RECT 258.305 128.345 258.535 130.100 ;
        RECT 258.785 128.345 259.015 130.100 ;
        RECT 259.225 130.075 259.500 130.100 ;
        RECT 259.225 128.350 259.550 130.075 ;
        RECT 259.265 128.345 259.495 128.350 ;
        RECT 259.745 128.345 259.975 130.100 ;
        RECT 260.225 129.525 260.455 131.345 ;
        RECT 260.705 131.275 260.935 131.345 ;
        RECT 260.650 130.100 260.975 131.275 ;
        RECT 260.175 128.350 260.500 129.525 ;
        RECT 260.225 128.345 260.455 128.350 ;
        RECT 260.705 128.345 260.935 130.100 ;
        RECT 261.185 129.525 261.415 131.345 ;
        RECT 261.665 131.275 261.895 131.345 ;
        RECT 261.625 130.100 261.950 131.275 ;
        RECT 261.125 128.350 261.475 129.525 ;
        RECT 261.185 128.345 261.415 128.350 ;
        RECT 261.665 128.345 261.895 130.100 ;
        RECT 262.145 129.525 262.375 131.345 ;
        RECT 262.625 131.275 262.855 131.345 ;
        RECT 262.575 130.100 262.900 131.275 ;
        RECT 262.100 128.350 262.425 129.525 ;
        RECT 262.145 128.345 262.375 128.350 ;
        RECT 262.625 128.345 262.855 130.100 ;
        RECT 263.105 129.525 263.335 131.345 ;
        RECT 263.585 131.275 263.815 131.345 ;
        RECT 263.525 130.100 263.875 131.275 ;
        RECT 263.050 128.350 263.375 129.525 ;
        RECT 263.105 128.345 263.335 128.350 ;
        RECT 263.585 128.345 263.815 130.100 ;
        RECT 264.065 129.525 264.295 131.345 ;
        RECT 264.545 131.275 264.775 131.345 ;
        RECT 264.500 130.100 264.825 131.275 ;
        RECT 264.025 128.350 264.350 129.525 ;
        RECT 264.065 128.345 264.295 128.350 ;
        RECT 264.545 128.345 264.775 130.100 ;
        RECT 265.025 129.525 265.255 131.345 ;
        RECT 265.505 131.275 265.735 131.345 ;
        RECT 265.450 130.100 265.775 131.275 ;
        RECT 264.975 128.350 265.300 129.525 ;
        RECT 265.025 128.345 265.255 128.350 ;
        RECT 265.505 128.345 265.735 130.100 ;
        RECT 265.985 129.525 266.215 131.345 ;
        RECT 266.465 131.275 266.695 131.345 ;
        RECT 266.425 130.100 266.750 131.275 ;
        RECT 265.925 128.350 266.250 129.525 ;
        RECT 265.985 128.345 266.215 128.350 ;
        RECT 266.465 128.345 266.695 130.100 ;
        RECT 266.945 129.525 267.175 131.345 ;
        RECT 267.425 131.275 267.655 131.345 ;
        RECT 267.375 130.100 267.700 131.275 ;
        RECT 266.900 128.350 267.225 129.525 ;
        RECT 266.945 128.345 267.175 128.350 ;
        RECT 267.425 128.345 267.655 130.100 ;
        RECT 267.905 129.525 268.135 131.345 ;
        RECT 268.385 131.275 268.615 131.345 ;
        RECT 268.865 131.275 269.095 131.345 ;
        RECT 269.345 131.275 269.575 131.345 ;
        RECT 269.825 131.275 270.055 131.345 ;
        RECT 270.305 131.275 270.535 131.345 ;
        RECT 268.325 130.100 270.575 131.275 ;
        RECT 267.850 128.350 268.175 129.525 ;
        RECT 267.905 128.345 268.135 128.350 ;
        RECT 268.385 128.345 268.615 130.100 ;
        RECT 268.865 128.345 269.095 130.100 ;
        RECT 269.345 128.345 269.575 130.100 ;
        RECT 269.825 128.345 270.055 130.100 ;
        RECT 270.305 128.345 270.535 130.100 ;
        RECT 257.525 126.150 270.350 128.150 ;
        RECT 257.345 125.300 257.575 125.950 ;
        RECT 257.825 125.300 258.055 125.950 ;
        RECT 258.305 125.300 258.535 125.950 ;
        RECT 258.785 125.300 259.015 125.950 ;
        RECT 259.225 125.325 259.550 125.950 ;
        RECT 259.225 125.300 259.525 125.325 ;
        RECT 259.745 125.300 259.975 125.950 ;
        RECT 260.175 125.550 260.500 125.950 ;
        RECT 257.300 124.900 259.525 125.300 ;
        RECT 259.700 124.900 260.025 125.300 ;
        RECT 260.225 124.950 260.455 125.550 ;
        RECT 260.705 125.300 260.935 125.950 ;
        RECT 261.125 125.550 261.475 125.950 ;
        RECT 260.650 124.900 261.000 125.300 ;
        RECT 261.185 124.950 261.415 125.550 ;
        RECT 261.665 125.300 261.895 125.950 ;
        RECT 262.100 125.550 262.425 125.950 ;
        RECT 261.625 124.900 261.950 125.300 ;
        RECT 262.145 124.950 262.375 125.550 ;
        RECT 262.625 125.300 262.855 125.950 ;
        RECT 263.050 125.550 263.375 125.950 ;
        RECT 262.575 124.900 262.900 125.300 ;
        RECT 263.105 124.950 263.335 125.550 ;
        RECT 263.585 125.300 263.815 125.950 ;
        RECT 264.025 125.550 264.350 125.950 ;
        RECT 263.525 124.900 263.875 125.300 ;
        RECT 264.065 124.950 264.295 125.550 ;
        RECT 264.545 125.300 264.775 125.950 ;
        RECT 264.975 125.550 265.300 125.950 ;
        RECT 264.500 124.900 264.825 125.300 ;
        RECT 265.025 124.950 265.255 125.550 ;
        RECT 265.505 125.300 265.735 125.950 ;
        RECT 265.925 125.550 266.275 125.950 ;
        RECT 265.450 124.900 265.800 125.300 ;
        RECT 265.985 124.950 266.215 125.550 ;
        RECT 266.465 125.300 266.695 125.950 ;
        RECT 266.900 125.550 267.225 125.950 ;
        RECT 266.425 124.900 266.750 125.300 ;
        RECT 266.945 124.950 267.175 125.550 ;
        RECT 267.425 125.300 267.655 125.950 ;
        RECT 267.850 125.550 268.200 125.950 ;
        RECT 267.375 124.900 267.700 125.300 ;
        RECT 267.905 124.950 268.135 125.550 ;
        RECT 268.385 125.300 268.615 125.950 ;
        RECT 268.865 125.300 269.095 125.950 ;
        RECT 269.345 125.300 269.575 125.950 ;
        RECT 269.825 125.300 270.055 125.950 ;
        RECT 270.305 125.300 270.535 125.950 ;
        RECT 268.325 124.900 270.575 125.300 ;
        RECT 270.900 124.750 271.250 131.550 ;
        RECT 236.370 124.745 236.600 124.750 ;
        RECT 236.850 124.745 237.080 124.750 ;
        RECT 237.330 124.745 237.560 124.750 ;
        RECT 237.810 124.745 238.040 124.750 ;
        RECT 238.290 124.745 238.520 124.750 ;
        RECT 240.970 124.745 241.200 124.750 ;
        RECT 241.450 124.745 241.680 124.750 ;
        RECT 241.930 124.745 242.160 124.750 ;
        RECT 242.410 124.745 242.640 124.750 ;
        RECT 242.890 124.745 243.120 124.750 ;
        RECT 245.570 124.745 245.800 124.750 ;
        RECT 246.050 124.745 246.280 124.750 ;
        RECT 246.530 124.745 246.760 124.750 ;
        RECT 247.010 124.745 247.240 124.750 ;
        RECT 247.490 124.745 247.720 124.750 ;
        RECT 237.050 124.545 237.850 124.550 ;
        RECT 242.100 124.545 242.475 124.550 ;
        RECT 246.250 124.545 247.050 124.550 ;
        RECT 230.000 123.225 232.975 123.825 ;
        RECT 129.370 122.035 129.620 122.075 ;
        RECT 130.200 122.035 130.450 122.075 ;
        RECT 131.030 122.035 131.280 122.075 ;
        RECT 131.860 122.035 132.110 122.075 ;
        RECT 132.690 122.035 132.940 122.075 ;
        RECT 133.520 122.035 133.770 122.075 ;
        RECT 134.350 122.035 134.600 122.075 ;
        RECT 135.180 122.035 135.430 122.075 ;
        RECT 136.010 122.035 136.260 122.075 ;
        RECT 136.840 122.035 137.090 122.075 ;
        RECT 137.670 122.035 137.920 122.075 ;
        RECT 138.500 122.035 138.750 122.075 ;
        RECT 139.330 122.035 139.580 122.075 ;
        RECT 140.160 122.035 140.410 122.075 ;
        RECT 140.990 122.035 141.240 122.075 ;
        RECT 141.820 122.035 142.070 122.075 ;
        RECT 142.650 122.035 142.900 122.075 ;
        RECT 143.480 122.035 143.730 122.075 ;
        RECT 144.310 122.035 144.560 122.075 ;
        RECT 145.140 122.035 145.390 122.075 ;
        RECT 145.970 122.035 146.220 122.075 ;
        RECT 146.800 122.035 147.050 122.075 ;
        RECT 147.630 122.035 147.880 122.075 ;
        RECT 148.460 122.035 148.710 122.075 ;
        RECT 149.290 122.035 149.540 122.075 ;
        RECT 150.120 122.035 150.370 122.075 ;
        RECT 150.950 122.035 151.200 122.075 ;
        RECT 151.780 122.035 152.030 122.075 ;
        RECT 152.610 122.035 152.860 122.075 ;
        RECT 153.440 122.035 153.690 122.075 ;
        RECT 154.270 122.035 154.520 122.075 ;
        RECT 155.100 122.035 155.350 122.075 ;
        RECT 155.930 122.035 156.180 122.075 ;
        RECT 156.760 122.035 157.010 122.075 ;
        RECT 157.590 122.035 157.840 122.075 ;
        RECT 158.420 122.035 158.670 122.075 ;
        RECT 159.250 122.035 159.500 122.075 ;
        RECT 160.080 122.035 160.330 122.075 ;
        RECT 160.910 122.035 161.160 122.075 ;
        RECT 161.740 122.035 161.990 122.075 ;
        RECT 162.570 122.035 162.820 122.075 ;
        RECT 163.400 122.035 163.650 122.075 ;
        RECT 164.230 122.035 164.480 122.075 ;
        RECT 165.060 122.035 165.310 122.075 ;
        RECT 165.890 122.035 166.140 122.075 ;
        RECT 166.720 122.035 166.970 122.075 ;
        RECT 167.550 122.035 167.800 122.075 ;
        RECT 168.380 122.035 168.630 122.075 ;
        RECT 169.210 122.035 169.460 122.075 ;
        RECT 170.040 122.035 170.290 122.075 ;
        RECT 170.870 122.035 171.120 122.075 ;
        RECT 171.700 122.035 171.950 122.075 ;
        RECT 172.530 122.035 172.780 122.075 ;
        RECT 173.360 122.035 173.610 122.075 ;
        RECT 174.190 122.035 174.440 122.075 ;
        RECT 175.020 122.035 175.270 122.075 ;
        RECT 175.850 122.035 176.100 122.075 ;
        RECT 176.680 122.035 176.930 122.075 ;
        RECT 177.510 122.035 177.760 122.075 ;
        RECT 178.340 122.035 178.590 122.075 ;
        RECT 179.170 122.035 179.420 122.075 ;
        RECT 180.000 122.035 180.250 122.075 ;
        RECT 180.830 122.035 181.080 122.075 ;
        RECT 181.660 122.035 181.910 122.075 ;
        RECT 182.490 122.035 182.740 122.075 ;
        RECT 183.320 122.035 183.570 122.075 ;
        RECT 184.150 122.035 184.400 122.075 ;
        RECT 184.980 122.035 185.230 122.075 ;
        RECT 185.810 122.035 186.060 122.075 ;
        RECT 186.640 122.035 186.890 122.075 ;
        RECT 187.470 122.035 187.720 122.075 ;
        RECT 188.300 122.035 188.550 122.075 ;
        RECT 189.130 122.035 189.380 122.075 ;
        RECT 189.960 122.035 190.210 122.075 ;
        RECT 190.790 122.035 191.040 122.075 ;
        RECT 191.620 122.035 191.870 122.075 ;
        RECT 192.450 122.035 192.700 122.075 ;
        RECT 193.280 122.035 193.530 122.075 ;
        RECT 194.110 122.035 194.360 122.075 ;
        RECT 194.940 122.035 195.190 122.075 ;
        RECT 195.770 122.035 196.020 122.075 ;
        RECT 196.600 122.035 196.850 122.075 ;
        RECT 197.430 122.035 197.680 122.075 ;
        RECT 198.260 122.035 198.510 122.075 ;
        RECT 199.090 122.035 199.340 122.075 ;
        RECT 199.920 122.035 200.170 122.075 ;
        RECT 200.750 122.035 201.000 122.075 ;
        RECT 201.580 122.035 201.830 122.075 ;
        RECT 202.410 122.035 202.660 122.075 ;
        RECT 203.240 122.035 203.490 122.075 ;
        RECT 204.070 122.035 204.320 122.075 ;
        RECT 204.900 122.035 205.150 122.075 ;
        RECT 205.730 122.035 205.980 122.075 ;
        RECT 206.560 122.035 206.810 122.075 ;
        RECT 207.390 122.035 207.640 122.075 ;
        RECT 208.220 122.035 208.470 122.075 ;
        RECT 209.050 122.035 209.300 122.075 ;
        RECT 209.880 122.035 210.130 122.075 ;
        RECT 210.710 122.035 210.960 122.075 ;
        RECT 211.540 122.035 211.790 122.075 ;
        RECT 212.325 121.525 231.425 122.350 ;
        RECT 75.275 120.650 231.425 121.525 ;
        RECT 231.775 121.350 232.025 123.225 ;
        RECT 232.200 121.350 232.550 122.350 ;
        RECT 232.725 121.350 232.975 123.225 ;
        RECT 233.325 122.350 233.700 124.500 ;
        RECT 237.045 124.170 237.850 124.545 ;
        RECT 242.095 124.170 242.475 124.545 ;
        RECT 246.245 124.170 247.050 124.545 ;
        RECT 237.050 123.825 237.850 124.170 ;
        RECT 242.100 123.825 242.475 124.170 ;
        RECT 246.250 123.825 247.050 124.170 ;
        RECT 250.825 124.175 253.580 124.550 ;
        RECT 256.625 124.425 271.250 124.750 ;
        RECT 250.825 123.825 253.575 124.175 ;
        RECT 256.625 123.900 271.250 124.250 ;
        RECT 234.900 123.225 237.850 123.825 ;
        RECT 239.500 123.225 242.475 123.825 ;
        RECT 244.775 123.225 247.050 123.825 ;
        RECT 248.700 123.225 253.575 123.825 ;
        RECT 237.050 122.550 237.850 123.225 ;
        RECT 242.100 122.550 242.475 123.225 ;
        RECT 246.250 122.550 247.050 123.225 ;
        RECT 250.825 122.875 253.575 123.225 ;
        RECT 250.825 122.550 253.580 122.875 ;
        RECT 233.325 121.350 237.085 122.350 ;
        RECT 237.275 121.350 237.625 122.350 ;
        RECT 237.815 121.350 239.250 122.350 ;
        RECT 231.950 120.825 232.800 121.150 ;
        RECT 233.325 120.650 236.650 121.350 ;
        RECT 238.250 120.650 239.250 121.350 ;
        RECT 240.250 121.350 241.685 122.350 ;
        RECT 241.875 121.350 242.225 122.350 ;
        RECT 242.415 121.350 243.850 122.350 ;
        RECT 240.250 121.150 241.250 121.350 ;
        RECT 242.850 121.150 243.850 121.350 ;
        RECT 240.250 120.650 241.525 121.150 ;
        RECT 242.575 120.650 243.850 121.150 ;
        RECT 244.850 121.350 246.285 122.350 ;
        RECT 246.475 121.350 246.825 122.350 ;
        RECT 247.015 121.350 250.880 122.350 ;
        RECT 251.075 121.350 251.400 122.350 ;
        RECT 244.850 120.650 245.850 121.350 ;
        RECT 247.450 121.325 250.880 121.350 ;
        RECT 247.450 120.650 250.875 121.325 ;
        RECT 251.600 120.650 251.850 122.350 ;
        RECT 252.050 121.350 252.375 122.350 ;
        RECT 252.550 120.650 252.800 122.350 ;
        RECT 253.000 121.350 253.325 122.350 ;
        RECT 253.525 120.800 254.950 122.350 ;
        RECT 253.525 120.650 263.775 120.800 ;
        RECT 75.275 119.450 263.775 120.650 ;
        RECT 75.275 110.200 228.050 119.450 ;
        RECT 272.800 114.675 273.400 166.450 ;
        RECT 56.450 104.375 228.050 110.200 ;
        RECT 56.450 104.275 97.300 104.375 ;
        RECT 75.275 100.500 97.300 104.275 ;
        RECT 97.830 103.825 98.080 103.860 ;
        RECT 98.660 103.825 98.910 103.860 ;
        RECT 99.490 103.825 99.740 103.860 ;
        RECT 100.320 103.825 100.570 103.860 ;
        RECT 101.150 103.825 101.400 103.860 ;
        RECT 101.980 103.825 102.230 103.860 ;
        RECT 102.810 103.825 103.060 103.860 ;
        RECT 103.640 103.825 103.890 103.860 ;
        RECT 104.470 103.825 104.720 103.860 ;
        RECT 105.300 103.825 105.550 103.860 ;
        RECT 106.130 103.825 106.380 103.860 ;
        RECT 106.960 103.825 107.210 103.860 ;
        RECT 107.790 103.825 108.040 103.860 ;
        RECT 108.620 103.825 108.870 103.860 ;
        RECT 109.450 103.825 109.700 103.860 ;
        RECT 110.280 103.825 110.530 103.860 ;
        RECT 111.110 103.825 111.360 103.860 ;
        RECT 111.940 103.825 112.190 103.860 ;
        RECT 112.770 103.825 113.020 103.860 ;
        RECT 113.600 103.825 113.850 103.860 ;
        RECT 114.430 103.825 114.680 103.860 ;
        RECT 115.260 103.825 115.510 103.860 ;
        RECT 116.090 103.825 116.340 103.860 ;
        RECT 116.920 103.825 117.170 103.860 ;
        RECT 117.750 103.825 118.000 103.860 ;
        RECT 118.580 103.825 118.830 103.860 ;
        RECT 119.410 103.825 119.660 103.860 ;
        RECT 120.240 103.825 120.490 103.860 ;
        RECT 121.070 103.825 121.320 103.860 ;
        RECT 121.900 103.825 122.150 103.860 ;
        RECT 122.730 103.825 122.980 103.860 ;
        RECT 123.560 103.825 123.810 103.860 ;
        RECT 124.390 103.825 124.640 103.860 ;
        RECT 125.220 103.825 125.470 103.860 ;
        RECT 126.050 103.825 126.300 103.860 ;
        RECT 126.880 103.825 127.130 103.860 ;
        RECT 97.825 101.800 98.925 103.825 ;
        RECT 99.475 101.800 100.575 103.825 ;
        RECT 101.150 101.800 102.250 103.825 ;
        RECT 102.800 101.800 103.900 103.825 ;
        RECT 104.470 101.800 105.575 103.825 ;
        RECT 106.125 101.800 107.225 103.825 ;
        RECT 107.790 101.800 108.900 103.825 ;
        RECT 109.450 101.800 110.550 103.825 ;
        RECT 111.100 101.800 112.200 103.825 ;
        RECT 112.770 101.800 113.875 103.825 ;
        RECT 114.425 101.800 115.525 103.825 ;
        RECT 116.090 101.800 117.200 103.825 ;
        RECT 117.750 101.800 118.850 103.825 ;
        RECT 119.400 101.800 120.500 103.825 ;
        RECT 121.070 101.800 122.175 103.825 ;
        RECT 122.725 101.800 123.825 103.825 ;
        RECT 124.390 101.800 125.500 103.825 ;
        RECT 126.050 101.800 127.150 103.825 ;
        RECT 97.830 101.755 98.080 101.800 ;
        RECT 98.660 101.755 98.910 101.800 ;
        RECT 99.490 101.755 99.740 101.800 ;
        RECT 100.320 101.755 100.570 101.800 ;
        RECT 101.150 101.755 101.400 101.800 ;
        RECT 101.980 101.755 102.230 101.800 ;
        RECT 102.810 101.755 103.060 101.800 ;
        RECT 103.640 101.755 103.890 101.800 ;
        RECT 104.470 101.755 104.720 101.800 ;
        RECT 105.300 101.755 105.550 101.800 ;
        RECT 106.130 101.755 106.380 101.800 ;
        RECT 106.960 101.755 107.210 101.800 ;
        RECT 107.790 101.755 108.040 101.800 ;
        RECT 108.620 101.755 108.870 101.800 ;
        RECT 109.450 101.755 109.700 101.800 ;
        RECT 110.280 101.755 110.530 101.800 ;
        RECT 111.110 101.755 111.360 101.800 ;
        RECT 111.940 101.755 112.190 101.800 ;
        RECT 112.770 101.755 113.020 101.800 ;
        RECT 113.600 101.755 113.850 101.800 ;
        RECT 114.430 101.755 114.680 101.800 ;
        RECT 115.260 101.755 115.510 101.800 ;
        RECT 116.090 101.755 116.340 101.800 ;
        RECT 116.920 101.755 117.170 101.800 ;
        RECT 117.750 101.755 118.000 101.800 ;
        RECT 118.580 101.755 118.830 101.800 ;
        RECT 119.410 101.755 119.660 101.800 ;
        RECT 120.240 101.755 120.490 101.800 ;
        RECT 121.070 101.755 121.320 101.800 ;
        RECT 121.900 101.755 122.150 101.800 ;
        RECT 122.730 101.755 122.980 101.800 ;
        RECT 123.560 101.755 123.810 101.800 ;
        RECT 124.390 101.755 124.640 101.800 ;
        RECT 125.220 101.755 125.470 101.800 ;
        RECT 126.050 101.755 126.300 101.800 ;
        RECT 126.880 101.755 127.130 101.800 ;
        RECT 127.675 101.750 128.825 103.875 ;
        RECT 129.370 103.825 129.620 103.860 ;
        RECT 130.200 103.825 130.450 103.860 ;
        RECT 131.030 103.825 131.280 103.860 ;
        RECT 131.860 103.825 132.110 103.860 ;
        RECT 132.690 103.825 132.940 103.860 ;
        RECT 133.520 103.825 133.770 103.860 ;
        RECT 134.350 103.825 134.600 103.860 ;
        RECT 135.180 103.825 135.430 103.860 ;
        RECT 136.010 103.825 136.260 103.860 ;
        RECT 136.840 103.825 137.090 103.860 ;
        RECT 137.670 103.825 137.920 103.860 ;
        RECT 138.500 103.825 138.750 103.860 ;
        RECT 139.330 103.825 139.580 103.860 ;
        RECT 140.160 103.825 140.410 103.860 ;
        RECT 140.990 103.825 141.240 103.860 ;
        RECT 141.820 103.825 142.070 103.860 ;
        RECT 142.650 103.825 142.900 103.860 ;
        RECT 143.480 103.825 143.730 103.860 ;
        RECT 144.310 103.825 144.560 103.860 ;
        RECT 145.140 103.825 145.390 103.860 ;
        RECT 145.970 103.825 146.220 103.860 ;
        RECT 146.800 103.825 147.050 103.860 ;
        RECT 147.630 103.825 147.880 103.860 ;
        RECT 148.460 103.825 148.710 103.860 ;
        RECT 149.290 103.825 149.540 103.860 ;
        RECT 150.120 103.825 150.370 103.860 ;
        RECT 150.950 103.825 151.200 103.860 ;
        RECT 151.780 103.825 152.030 103.860 ;
        RECT 152.610 103.825 152.860 103.860 ;
        RECT 153.440 103.825 153.690 103.860 ;
        RECT 154.270 103.825 154.520 103.860 ;
        RECT 155.100 103.825 155.350 103.860 ;
        RECT 155.930 103.825 156.180 103.860 ;
        RECT 156.760 103.825 157.010 103.860 ;
        RECT 157.590 103.825 157.840 103.860 ;
        RECT 158.420 103.825 158.670 103.860 ;
        RECT 159.250 103.825 159.500 103.860 ;
        RECT 160.080 103.825 160.330 103.860 ;
        RECT 160.910 103.825 161.160 103.860 ;
        RECT 161.740 103.825 161.990 103.860 ;
        RECT 162.570 103.825 162.820 103.860 ;
        RECT 163.400 103.825 163.650 103.860 ;
        RECT 164.230 103.825 164.480 103.860 ;
        RECT 165.060 103.825 165.310 103.860 ;
        RECT 165.890 103.825 166.140 103.860 ;
        RECT 166.720 103.825 166.970 103.860 ;
        RECT 167.550 103.825 167.800 103.860 ;
        RECT 168.380 103.825 168.630 103.860 ;
        RECT 169.210 103.825 169.460 103.860 ;
        RECT 170.040 103.825 170.290 103.860 ;
        RECT 170.870 103.825 171.120 103.860 ;
        RECT 171.700 103.825 171.950 103.860 ;
        RECT 172.530 103.825 172.780 103.860 ;
        RECT 173.360 103.825 173.610 103.860 ;
        RECT 174.190 103.825 174.440 103.860 ;
        RECT 175.020 103.825 175.270 103.860 ;
        RECT 175.850 103.825 176.100 103.860 ;
        RECT 176.680 103.825 176.930 103.860 ;
        RECT 177.510 103.825 177.760 103.860 ;
        RECT 178.340 103.825 178.590 103.860 ;
        RECT 179.170 103.825 179.420 103.860 ;
        RECT 180.000 103.825 180.250 103.860 ;
        RECT 180.830 103.825 181.080 103.860 ;
        RECT 181.660 103.825 181.910 103.860 ;
        RECT 182.490 103.825 182.740 103.860 ;
        RECT 183.320 103.825 183.570 103.860 ;
        RECT 184.150 103.825 184.400 103.860 ;
        RECT 184.980 103.825 185.230 103.860 ;
        RECT 185.810 103.825 186.060 103.860 ;
        RECT 186.640 103.825 186.890 103.860 ;
        RECT 187.470 103.825 187.720 103.860 ;
        RECT 188.300 103.825 188.550 103.860 ;
        RECT 189.130 103.825 189.380 103.860 ;
        RECT 189.960 103.825 190.210 103.860 ;
        RECT 190.790 103.825 191.040 103.860 ;
        RECT 191.620 103.825 191.870 103.860 ;
        RECT 192.450 103.825 192.700 103.860 ;
        RECT 193.280 103.825 193.530 103.860 ;
        RECT 194.110 103.825 194.360 103.860 ;
        RECT 194.940 103.825 195.190 103.860 ;
        RECT 195.770 103.825 196.020 103.860 ;
        RECT 196.600 103.825 196.850 103.860 ;
        RECT 197.430 103.825 197.680 103.860 ;
        RECT 198.260 103.825 198.510 103.860 ;
        RECT 199.090 103.825 199.340 103.860 ;
        RECT 199.920 103.825 200.170 103.860 ;
        RECT 200.750 103.825 201.000 103.860 ;
        RECT 201.580 103.825 201.830 103.860 ;
        RECT 202.410 103.825 202.660 103.860 ;
        RECT 203.240 103.825 203.490 103.860 ;
        RECT 204.070 103.825 204.320 103.860 ;
        RECT 204.900 103.825 205.150 103.860 ;
        RECT 205.730 103.825 205.980 103.860 ;
        RECT 206.560 103.825 206.810 103.860 ;
        RECT 207.390 103.825 207.640 103.860 ;
        RECT 208.220 103.825 208.470 103.860 ;
        RECT 209.050 103.825 209.300 103.860 ;
        RECT 209.880 103.825 210.130 103.860 ;
        RECT 210.710 103.825 210.960 103.860 ;
        RECT 211.540 103.825 211.790 103.860 ;
        RECT 129.370 101.800 130.475 103.825 ;
        RECT 131.025 101.800 132.125 103.825 ;
        RECT 132.690 101.800 133.800 103.825 ;
        RECT 134.350 101.800 135.450 103.825 ;
        RECT 136.000 101.800 137.100 103.825 ;
        RECT 137.670 101.800 138.775 103.825 ;
        RECT 139.325 101.800 140.425 103.825 ;
        RECT 140.990 101.800 142.100 103.825 ;
        RECT 142.650 101.800 143.750 103.825 ;
        RECT 144.300 101.800 145.400 103.825 ;
        RECT 145.950 101.800 147.050 103.825 ;
        RECT 147.625 101.800 148.725 103.825 ;
        RECT 149.290 101.800 150.400 103.825 ;
        RECT 150.950 101.800 152.050 103.825 ;
        RECT 152.600 101.800 153.700 103.825 ;
        RECT 154.270 101.800 155.375 103.825 ;
        RECT 155.925 101.800 157.025 103.825 ;
        RECT 157.575 101.800 158.675 103.825 ;
        RECT 159.250 101.800 160.350 103.825 ;
        RECT 160.900 101.800 162.000 103.825 ;
        RECT 162.570 101.800 163.675 103.825 ;
        RECT 164.225 101.800 165.325 103.825 ;
        RECT 165.890 101.800 167.000 103.825 ;
        RECT 167.550 101.800 168.650 103.825 ;
        RECT 169.200 101.800 170.300 103.825 ;
        RECT 170.870 101.800 171.975 103.825 ;
        RECT 172.525 101.800 173.625 103.825 ;
        RECT 174.190 101.800 175.300 103.825 ;
        RECT 175.850 101.800 176.950 103.825 ;
        RECT 177.500 101.800 178.600 103.825 ;
        RECT 179.170 101.800 180.275 103.825 ;
        RECT 180.825 101.800 181.925 103.825 ;
        RECT 182.490 101.800 183.600 103.825 ;
        RECT 184.150 101.800 185.250 103.825 ;
        RECT 185.800 101.800 186.900 103.825 ;
        RECT 187.470 101.800 188.575 103.825 ;
        RECT 189.125 101.800 190.225 103.825 ;
        RECT 190.790 101.800 191.900 103.825 ;
        RECT 192.450 101.800 193.550 103.825 ;
        RECT 194.100 101.800 195.200 103.825 ;
        RECT 195.770 101.800 196.875 103.825 ;
        RECT 197.425 101.800 198.525 103.825 ;
        RECT 199.090 101.800 200.200 103.825 ;
        RECT 200.750 101.800 201.850 103.825 ;
        RECT 202.400 101.800 203.500 103.825 ;
        RECT 204.070 101.800 205.175 103.825 ;
        RECT 205.725 101.800 206.825 103.825 ;
        RECT 207.390 101.800 208.500 103.825 ;
        RECT 209.050 101.800 210.150 103.825 ;
        RECT 210.700 101.800 211.800 103.825 ;
        RECT 129.370 101.755 129.620 101.800 ;
        RECT 130.200 101.755 130.450 101.800 ;
        RECT 131.030 101.755 131.280 101.800 ;
        RECT 131.860 101.755 132.110 101.800 ;
        RECT 132.690 101.755 132.940 101.800 ;
        RECT 133.520 101.755 133.770 101.800 ;
        RECT 134.350 101.755 134.600 101.800 ;
        RECT 135.180 101.755 135.430 101.800 ;
        RECT 136.010 101.755 136.260 101.800 ;
        RECT 136.840 101.755 137.090 101.800 ;
        RECT 137.670 101.755 137.920 101.800 ;
        RECT 138.500 101.755 138.750 101.800 ;
        RECT 139.330 101.755 139.580 101.800 ;
        RECT 140.160 101.755 140.410 101.800 ;
        RECT 140.990 101.755 141.240 101.800 ;
        RECT 141.820 101.755 142.070 101.800 ;
        RECT 142.650 101.755 142.900 101.800 ;
        RECT 143.480 101.755 143.730 101.800 ;
        RECT 144.310 101.755 144.560 101.800 ;
        RECT 145.140 101.755 145.390 101.800 ;
        RECT 145.970 101.755 146.220 101.800 ;
        RECT 146.800 101.755 147.050 101.800 ;
        RECT 147.630 101.755 147.880 101.800 ;
        RECT 148.460 101.755 148.710 101.800 ;
        RECT 149.290 101.755 149.540 101.800 ;
        RECT 150.120 101.755 150.370 101.800 ;
        RECT 150.950 101.755 151.200 101.800 ;
        RECT 151.780 101.755 152.030 101.800 ;
        RECT 152.610 101.755 152.860 101.800 ;
        RECT 153.440 101.755 153.690 101.800 ;
        RECT 154.270 101.755 154.520 101.800 ;
        RECT 155.100 101.755 155.350 101.800 ;
        RECT 155.930 101.755 156.180 101.800 ;
        RECT 156.760 101.755 157.010 101.800 ;
        RECT 157.590 101.755 157.840 101.800 ;
        RECT 158.420 101.755 158.670 101.800 ;
        RECT 159.250 101.755 159.500 101.800 ;
        RECT 160.080 101.755 160.330 101.800 ;
        RECT 160.910 101.755 161.160 101.800 ;
        RECT 161.740 101.755 161.990 101.800 ;
        RECT 162.570 101.755 162.820 101.800 ;
        RECT 163.400 101.755 163.650 101.800 ;
        RECT 164.230 101.755 164.480 101.800 ;
        RECT 165.060 101.755 165.310 101.800 ;
        RECT 165.890 101.755 166.140 101.800 ;
        RECT 166.720 101.755 166.970 101.800 ;
        RECT 167.550 101.755 167.800 101.800 ;
        RECT 168.380 101.755 168.630 101.800 ;
        RECT 169.210 101.755 169.460 101.800 ;
        RECT 170.040 101.755 170.290 101.800 ;
        RECT 170.870 101.755 171.120 101.800 ;
        RECT 171.700 101.755 171.950 101.800 ;
        RECT 172.530 101.755 172.780 101.800 ;
        RECT 173.360 101.755 173.610 101.800 ;
        RECT 174.190 101.755 174.440 101.800 ;
        RECT 175.020 101.755 175.270 101.800 ;
        RECT 175.850 101.755 176.100 101.800 ;
        RECT 176.680 101.755 176.930 101.800 ;
        RECT 177.510 101.755 177.760 101.800 ;
        RECT 178.340 101.755 178.590 101.800 ;
        RECT 179.170 101.755 179.420 101.800 ;
        RECT 180.000 101.755 180.250 101.800 ;
        RECT 180.830 101.755 181.080 101.800 ;
        RECT 181.660 101.755 181.910 101.800 ;
        RECT 182.490 101.755 182.740 101.800 ;
        RECT 183.320 101.755 183.570 101.800 ;
        RECT 184.150 101.755 184.400 101.800 ;
        RECT 184.980 101.755 185.230 101.800 ;
        RECT 185.810 101.755 186.060 101.800 ;
        RECT 186.640 101.755 186.890 101.800 ;
        RECT 187.470 101.755 187.720 101.800 ;
        RECT 188.300 101.755 188.550 101.800 ;
        RECT 189.130 101.755 189.380 101.800 ;
        RECT 189.960 101.755 190.210 101.800 ;
        RECT 190.790 101.755 191.040 101.800 ;
        RECT 191.620 101.755 191.870 101.800 ;
        RECT 192.450 101.755 192.700 101.800 ;
        RECT 193.280 101.755 193.530 101.800 ;
        RECT 194.110 101.755 194.360 101.800 ;
        RECT 194.940 101.755 195.190 101.800 ;
        RECT 195.770 101.755 196.020 101.800 ;
        RECT 196.600 101.755 196.850 101.800 ;
        RECT 197.430 101.755 197.680 101.800 ;
        RECT 198.260 101.755 198.510 101.800 ;
        RECT 199.090 101.755 199.340 101.800 ;
        RECT 199.920 101.755 200.170 101.800 ;
        RECT 200.750 101.755 201.000 101.800 ;
        RECT 201.580 101.755 201.830 101.800 ;
        RECT 202.410 101.755 202.660 101.800 ;
        RECT 203.240 101.755 203.490 101.800 ;
        RECT 204.070 101.755 204.320 101.800 ;
        RECT 204.900 101.755 205.150 101.800 ;
        RECT 205.730 101.755 205.980 101.800 ;
        RECT 206.560 101.755 206.810 101.800 ;
        RECT 207.390 101.755 207.640 101.800 ;
        RECT 208.220 101.755 208.470 101.800 ;
        RECT 209.050 101.755 209.300 101.800 ;
        RECT 209.880 101.755 210.130 101.800 ;
        RECT 210.710 101.755 210.960 101.800 ;
        RECT 211.540 101.755 211.790 101.800 ;
        RECT 212.325 100.500 228.050 104.375 ;
        RECT 97.830 99.825 98.080 99.865 ;
        RECT 98.660 99.825 98.910 99.865 ;
        RECT 99.490 99.825 99.740 99.865 ;
        RECT 100.320 99.825 100.570 99.865 ;
        RECT 101.150 99.825 101.400 99.865 ;
        RECT 101.980 99.825 102.230 99.865 ;
        RECT 102.810 99.825 103.060 99.865 ;
        RECT 103.640 99.825 103.890 99.865 ;
        RECT 104.470 99.825 104.720 99.865 ;
        RECT 105.300 99.825 105.550 99.865 ;
        RECT 106.130 99.825 106.380 99.865 ;
        RECT 106.960 99.825 107.210 99.865 ;
        RECT 107.790 99.825 108.040 99.865 ;
        RECT 108.620 99.825 108.870 99.865 ;
        RECT 109.450 99.825 109.700 99.865 ;
        RECT 110.280 99.825 110.530 99.865 ;
        RECT 111.110 99.825 111.360 99.865 ;
        RECT 111.940 99.825 112.190 99.865 ;
        RECT 112.770 99.825 113.020 99.865 ;
        RECT 113.600 99.825 113.850 99.865 ;
        RECT 114.430 99.825 114.680 99.865 ;
        RECT 115.260 99.825 115.510 99.865 ;
        RECT 116.090 99.825 116.340 99.865 ;
        RECT 116.920 99.825 117.170 99.865 ;
        RECT 117.750 99.825 118.000 99.865 ;
        RECT 118.580 99.825 118.830 99.865 ;
        RECT 119.410 99.825 119.660 99.865 ;
        RECT 120.240 99.825 120.490 99.865 ;
        RECT 121.070 99.825 121.320 99.865 ;
        RECT 121.900 99.825 122.150 99.865 ;
        RECT 122.730 99.825 122.980 99.865 ;
        RECT 123.560 99.825 123.810 99.865 ;
        RECT 124.390 99.825 124.640 99.865 ;
        RECT 125.220 99.825 125.470 99.865 ;
        RECT 126.050 99.825 126.300 99.865 ;
        RECT 126.880 99.825 127.130 99.865 ;
        RECT 127.710 99.825 127.960 99.865 ;
        RECT 128.540 99.825 128.790 99.865 ;
        RECT 129.370 99.825 129.620 99.865 ;
        RECT 130.200 99.825 130.450 99.865 ;
        RECT 131.030 99.825 131.280 99.865 ;
        RECT 131.860 99.825 132.110 99.865 ;
        RECT 132.690 99.825 132.940 99.865 ;
        RECT 133.520 99.825 133.770 99.865 ;
        RECT 134.350 99.825 134.600 99.865 ;
        RECT 135.180 99.825 135.430 99.865 ;
        RECT 136.010 99.825 136.260 99.865 ;
        RECT 136.840 99.825 137.090 99.865 ;
        RECT 137.670 99.825 137.920 99.865 ;
        RECT 138.500 99.825 138.750 99.865 ;
        RECT 139.330 99.825 139.580 99.865 ;
        RECT 140.160 99.825 140.410 99.865 ;
        RECT 140.990 99.825 141.240 99.865 ;
        RECT 141.820 99.825 142.070 99.865 ;
        RECT 142.650 99.825 142.900 99.865 ;
        RECT 143.480 99.825 143.730 99.865 ;
        RECT 144.310 99.825 144.560 99.865 ;
        RECT 145.140 99.825 145.390 99.865 ;
        RECT 145.970 99.825 146.220 99.865 ;
        RECT 146.800 99.825 147.050 99.865 ;
        RECT 147.630 99.825 147.880 99.865 ;
        RECT 148.460 99.825 148.710 99.865 ;
        RECT 149.290 99.825 149.540 99.865 ;
        RECT 150.120 99.825 150.370 99.865 ;
        RECT 150.950 99.825 151.200 99.865 ;
        RECT 151.780 99.825 152.030 99.865 ;
        RECT 152.610 99.825 152.860 99.865 ;
        RECT 153.440 99.825 153.690 99.865 ;
        RECT 154.270 99.825 154.520 99.865 ;
        RECT 155.100 99.825 155.350 99.865 ;
        RECT 155.930 99.825 156.180 99.865 ;
        RECT 156.760 99.825 157.010 99.865 ;
        RECT 157.590 99.825 157.840 99.865 ;
        RECT 158.420 99.825 158.670 99.865 ;
        RECT 159.250 99.825 159.500 99.865 ;
        RECT 160.080 99.825 160.330 99.865 ;
        RECT 160.910 99.825 161.160 99.865 ;
        RECT 161.740 99.825 161.990 99.865 ;
        RECT 162.570 99.825 162.820 99.865 ;
        RECT 163.400 99.825 163.650 99.865 ;
        RECT 164.230 99.825 164.480 99.865 ;
        RECT 165.060 99.825 165.310 99.865 ;
        RECT 165.890 99.825 166.140 99.865 ;
        RECT 166.720 99.825 166.970 99.865 ;
        RECT 167.550 99.825 167.800 99.865 ;
        RECT 168.380 99.825 168.630 99.865 ;
        RECT 169.210 99.825 169.460 99.865 ;
        RECT 170.040 99.825 170.290 99.865 ;
        RECT 170.870 99.825 171.120 99.865 ;
        RECT 171.700 99.825 171.950 99.865 ;
        RECT 172.530 99.825 172.780 99.865 ;
        RECT 173.360 99.825 173.610 99.865 ;
        RECT 174.190 99.825 174.440 99.865 ;
        RECT 175.020 99.825 175.270 99.865 ;
        RECT 175.850 99.825 176.100 99.865 ;
        RECT 176.680 99.825 176.930 99.865 ;
        RECT 177.510 99.825 177.760 99.865 ;
        RECT 178.340 99.825 178.590 99.865 ;
        RECT 179.170 99.825 179.420 99.865 ;
        RECT 56.450 97.800 98.100 99.825 ;
        RECT 98.650 97.800 99.750 99.825 ;
        RECT 100.300 97.800 101.425 99.825 ;
        RECT 101.975 97.800 103.075 99.825 ;
        RECT 103.625 97.800 104.725 99.825 ;
        RECT 105.300 97.800 106.400 99.825 ;
        RECT 106.950 97.800 108.050 99.825 ;
        RECT 108.600 97.800 109.700 99.825 ;
        RECT 110.275 97.800 111.375 99.825 ;
        RECT 56.450 18.125 58.475 97.800 ;
        RECT 97.830 97.760 98.080 97.800 ;
        RECT 98.660 97.760 98.910 97.800 ;
        RECT 99.490 97.760 99.740 97.800 ;
        RECT 100.320 97.760 100.570 97.800 ;
        RECT 101.150 97.760 101.400 97.800 ;
        RECT 101.980 97.760 102.230 97.800 ;
        RECT 102.810 97.760 103.060 97.800 ;
        RECT 103.640 97.760 103.890 97.800 ;
        RECT 104.470 97.760 104.720 97.800 ;
        RECT 105.300 97.760 105.550 97.800 ;
        RECT 106.130 97.760 106.380 97.800 ;
        RECT 106.960 97.760 107.210 97.800 ;
        RECT 107.790 97.760 108.040 97.800 ;
        RECT 108.620 97.760 108.870 97.800 ;
        RECT 109.450 97.760 109.700 97.800 ;
        RECT 110.280 97.760 110.530 97.800 ;
        RECT 111.110 97.760 111.360 97.800 ;
        RECT 111.925 97.625 113.050 99.825 ;
        RECT 113.600 97.800 114.700 99.825 ;
        RECT 115.250 97.800 116.350 99.825 ;
        RECT 116.920 97.800 118.025 99.825 ;
        RECT 118.575 97.800 119.675 99.825 ;
        RECT 120.225 97.800 121.325 99.825 ;
        RECT 121.900 97.800 123.000 99.825 ;
        RECT 123.550 97.800 124.650 99.825 ;
        RECT 125.220 97.800 126.325 99.825 ;
        RECT 126.875 97.800 127.975 99.825 ;
        RECT 128.525 97.800 129.625 99.825 ;
        RECT 130.200 97.800 131.300 99.825 ;
        RECT 131.850 97.800 132.950 99.825 ;
        RECT 133.520 97.800 134.625 99.825 ;
        RECT 135.175 97.800 136.275 99.825 ;
        RECT 136.825 97.800 137.925 99.825 ;
        RECT 138.500 97.800 139.600 99.825 ;
        RECT 140.150 97.800 141.250 99.825 ;
        RECT 141.820 97.800 142.925 99.825 ;
        RECT 143.475 97.800 144.575 99.825 ;
        RECT 145.140 97.800 146.250 99.825 ;
        RECT 146.800 97.800 147.900 99.825 ;
        RECT 148.450 97.800 149.550 99.825 ;
        RECT 150.120 97.800 151.225 99.825 ;
        RECT 151.775 97.800 152.875 99.825 ;
        RECT 153.440 97.800 154.550 99.825 ;
        RECT 155.100 97.800 156.200 99.825 ;
        RECT 156.750 97.800 157.850 99.825 ;
        RECT 158.420 97.800 159.525 99.825 ;
        RECT 160.075 97.800 161.175 99.825 ;
        RECT 161.725 97.800 162.825 99.825 ;
        RECT 163.400 97.800 164.500 99.825 ;
        RECT 165.050 97.800 166.150 99.825 ;
        RECT 166.720 97.800 167.825 99.825 ;
        RECT 168.375 97.800 169.475 99.825 ;
        RECT 170.025 97.800 171.125 99.825 ;
        RECT 171.675 97.800 172.780 99.825 ;
        RECT 173.350 97.800 174.450 99.825 ;
        RECT 175.020 97.800 176.125 99.825 ;
        RECT 176.675 97.800 177.775 99.825 ;
        RECT 178.325 97.800 179.425 99.825 ;
        RECT 113.600 97.760 113.850 97.800 ;
        RECT 114.430 97.760 114.680 97.800 ;
        RECT 115.260 97.760 115.510 97.800 ;
        RECT 116.090 97.760 116.340 97.800 ;
        RECT 116.920 97.760 117.170 97.800 ;
        RECT 117.750 97.760 118.000 97.800 ;
        RECT 118.580 97.760 118.830 97.800 ;
        RECT 119.410 97.760 119.660 97.800 ;
        RECT 120.240 97.760 120.490 97.800 ;
        RECT 121.070 97.760 121.320 97.800 ;
        RECT 121.900 97.760 122.150 97.800 ;
        RECT 122.730 97.760 122.980 97.800 ;
        RECT 123.560 97.760 123.810 97.800 ;
        RECT 124.390 97.760 124.640 97.800 ;
        RECT 125.220 97.760 125.470 97.800 ;
        RECT 126.050 97.760 126.300 97.800 ;
        RECT 126.880 97.760 127.130 97.800 ;
        RECT 127.710 97.760 127.960 97.800 ;
        RECT 128.540 97.760 128.790 97.800 ;
        RECT 129.370 97.760 129.620 97.800 ;
        RECT 130.200 97.760 130.450 97.800 ;
        RECT 131.030 97.760 131.280 97.800 ;
        RECT 131.860 97.760 132.110 97.800 ;
        RECT 132.690 97.760 132.940 97.800 ;
        RECT 133.520 97.760 133.770 97.800 ;
        RECT 134.350 97.760 134.600 97.800 ;
        RECT 135.180 97.760 135.430 97.800 ;
        RECT 136.010 97.760 136.260 97.800 ;
        RECT 136.840 97.760 137.090 97.800 ;
        RECT 137.670 97.760 137.920 97.800 ;
        RECT 138.500 97.760 138.750 97.800 ;
        RECT 139.330 97.760 139.580 97.800 ;
        RECT 140.160 97.760 140.410 97.800 ;
        RECT 140.990 97.760 141.240 97.800 ;
        RECT 141.820 97.760 142.070 97.800 ;
        RECT 142.650 97.760 142.900 97.800 ;
        RECT 143.480 97.760 143.730 97.800 ;
        RECT 144.310 97.760 144.560 97.800 ;
        RECT 145.140 97.760 145.390 97.800 ;
        RECT 145.970 97.760 146.220 97.800 ;
        RECT 146.800 97.760 147.050 97.800 ;
        RECT 147.630 97.760 147.880 97.800 ;
        RECT 148.460 97.760 148.710 97.800 ;
        RECT 149.290 97.760 149.540 97.800 ;
        RECT 150.120 97.760 150.370 97.800 ;
        RECT 150.950 97.760 151.200 97.800 ;
        RECT 151.780 97.760 152.030 97.800 ;
        RECT 152.610 97.760 152.860 97.800 ;
        RECT 153.440 97.760 153.690 97.800 ;
        RECT 154.270 97.760 154.520 97.800 ;
        RECT 155.100 97.760 155.350 97.800 ;
        RECT 155.930 97.760 156.180 97.800 ;
        RECT 156.760 97.760 157.010 97.800 ;
        RECT 157.590 97.760 157.840 97.800 ;
        RECT 158.420 97.760 158.670 97.800 ;
        RECT 159.250 97.760 159.500 97.800 ;
        RECT 160.080 97.760 160.330 97.800 ;
        RECT 160.910 97.760 161.160 97.800 ;
        RECT 161.740 97.760 161.990 97.800 ;
        RECT 162.570 97.760 162.820 97.800 ;
        RECT 163.400 97.760 163.650 97.800 ;
        RECT 164.230 97.760 164.480 97.800 ;
        RECT 165.060 97.760 165.310 97.800 ;
        RECT 165.890 97.760 166.140 97.800 ;
        RECT 166.720 97.760 166.970 97.800 ;
        RECT 167.550 97.760 167.800 97.800 ;
        RECT 168.380 97.760 168.630 97.800 ;
        RECT 169.210 97.760 169.460 97.800 ;
        RECT 170.040 97.760 170.290 97.800 ;
        RECT 170.870 97.760 171.120 97.800 ;
        RECT 171.700 97.760 171.950 97.800 ;
        RECT 172.530 97.760 172.780 97.800 ;
        RECT 173.360 97.760 173.610 97.800 ;
        RECT 174.190 97.760 174.440 97.800 ;
        RECT 175.020 97.760 175.270 97.800 ;
        RECT 175.850 97.760 176.100 97.800 ;
        RECT 176.680 97.760 176.930 97.800 ;
        RECT 177.510 97.760 177.760 97.800 ;
        RECT 178.340 97.760 178.590 97.800 ;
        RECT 179.170 97.760 179.420 97.800 ;
        RECT 179.900 97.750 180.350 99.875 ;
        RECT 180.650 97.750 181.250 99.875 ;
        RECT 181.660 99.825 181.910 99.865 ;
        RECT 182.490 99.825 182.740 99.865 ;
        RECT 183.320 99.825 183.570 99.865 ;
        RECT 184.150 99.825 184.400 99.865 ;
        RECT 184.980 99.825 185.230 99.865 ;
        RECT 185.810 99.825 186.060 99.865 ;
        RECT 186.640 99.825 186.890 99.865 ;
        RECT 187.470 99.825 187.720 99.865 ;
        RECT 188.300 99.825 188.550 99.865 ;
        RECT 189.130 99.825 189.380 99.865 ;
        RECT 189.960 99.825 190.210 99.865 ;
        RECT 190.790 99.825 191.040 99.865 ;
        RECT 191.620 99.825 191.870 99.865 ;
        RECT 192.450 99.825 192.700 99.865 ;
        RECT 193.280 99.825 193.530 99.865 ;
        RECT 194.110 99.825 194.360 99.865 ;
        RECT 194.940 99.825 195.190 99.865 ;
        RECT 195.770 99.825 196.020 99.865 ;
        RECT 196.600 99.825 196.850 99.865 ;
        RECT 197.430 99.825 197.680 99.865 ;
        RECT 198.260 99.825 198.510 99.865 ;
        RECT 199.090 99.825 199.340 99.865 ;
        RECT 199.920 99.825 200.170 99.865 ;
        RECT 200.750 99.825 201.000 99.865 ;
        RECT 201.580 99.825 201.830 99.865 ;
        RECT 202.410 99.825 202.660 99.865 ;
        RECT 203.240 99.825 203.490 99.865 ;
        RECT 204.070 99.825 204.320 99.865 ;
        RECT 204.900 99.825 205.150 99.865 ;
        RECT 205.730 99.825 205.980 99.865 ;
        RECT 206.560 99.825 206.810 99.865 ;
        RECT 207.390 99.825 207.640 99.865 ;
        RECT 208.220 99.825 208.470 99.865 ;
        RECT 209.050 99.825 209.300 99.865 ;
        RECT 209.880 99.825 210.130 99.865 ;
        RECT 210.710 99.825 210.960 99.865 ;
        RECT 211.540 99.825 211.790 99.865 ;
        RECT 181.650 97.800 182.750 99.825 ;
        RECT 183.320 97.800 184.425 99.825 ;
        RECT 184.975 97.800 186.075 99.825 ;
        RECT 186.640 97.800 187.750 99.825 ;
        RECT 188.300 97.800 189.400 99.825 ;
        RECT 189.950 97.800 191.050 99.825 ;
        RECT 191.600 97.800 192.700 99.825 ;
        RECT 193.275 97.800 194.375 99.825 ;
        RECT 194.925 97.800 196.025 99.825 ;
        RECT 196.575 97.800 197.680 99.825 ;
        RECT 198.250 97.800 199.350 99.825 ;
        RECT 199.920 97.800 201.025 99.825 ;
        RECT 201.575 97.800 202.675 99.825 ;
        RECT 203.225 97.800 204.325 99.825 ;
        RECT 204.900 97.800 206.000 99.825 ;
        RECT 206.550 97.800 207.650 99.825 ;
        RECT 208.200 97.800 209.300 99.825 ;
        RECT 209.875 97.800 210.975 99.825 ;
        RECT 211.525 97.800 214.125 99.825 ;
        RECT 181.660 97.760 181.910 97.800 ;
        RECT 182.490 97.760 182.740 97.800 ;
        RECT 183.320 97.760 183.570 97.800 ;
        RECT 184.150 97.760 184.400 97.800 ;
        RECT 184.980 97.760 185.230 97.800 ;
        RECT 185.810 97.760 186.060 97.800 ;
        RECT 186.640 97.760 186.890 97.800 ;
        RECT 187.470 97.760 187.720 97.800 ;
        RECT 188.300 97.760 188.550 97.800 ;
        RECT 189.130 97.760 189.380 97.800 ;
        RECT 189.960 97.760 190.210 97.800 ;
        RECT 190.790 97.760 191.040 97.800 ;
        RECT 191.620 97.760 191.870 97.800 ;
        RECT 192.450 97.760 192.700 97.800 ;
        RECT 193.280 97.760 193.530 97.800 ;
        RECT 194.110 97.760 194.360 97.800 ;
        RECT 194.940 97.760 195.190 97.800 ;
        RECT 195.770 97.760 196.020 97.800 ;
        RECT 196.600 97.760 196.850 97.800 ;
        RECT 197.430 97.760 197.680 97.800 ;
        RECT 198.260 97.760 198.510 97.800 ;
        RECT 199.090 97.760 199.340 97.800 ;
        RECT 199.920 97.760 200.170 97.800 ;
        RECT 200.750 97.760 201.000 97.800 ;
        RECT 201.580 97.760 201.830 97.800 ;
        RECT 202.410 97.760 202.660 97.800 ;
        RECT 203.240 97.760 203.490 97.800 ;
        RECT 204.070 97.760 204.320 97.800 ;
        RECT 204.900 97.760 205.150 97.800 ;
        RECT 205.730 97.760 205.980 97.800 ;
        RECT 206.560 97.760 206.810 97.800 ;
        RECT 207.390 97.760 207.640 97.800 ;
        RECT 208.220 97.760 208.470 97.800 ;
        RECT 209.050 97.760 209.300 97.800 ;
        RECT 209.880 97.760 210.130 97.800 ;
        RECT 210.710 97.760 210.960 97.800 ;
        RECT 211.540 97.760 211.790 97.800 ;
        RECT 215.625 97.100 228.050 100.500 ;
        RECT 65.000 96.395 75.900 96.400 ;
        RECT 65.000 95.645 226.130 96.395 ;
        RECT 65.000 94.675 84.705 95.645 ;
        RECT 75.280 93.595 84.705 94.675 ;
        RECT 75.280 84.295 77.805 93.595 ;
        RECT 78.305 84.295 79.105 93.320 ;
        RECT 79.580 84.295 80.380 93.595 ;
        RECT 80.855 84.295 81.655 93.320 ;
        RECT 82.155 84.295 84.705 93.595 ;
        RECT 86.030 95.620 98.030 95.645 ;
        RECT 86.030 93.320 86.780 95.620 ;
        RECT 87.030 93.750 87.880 95.170 ;
        RECT 88.230 94.820 95.805 95.620 ;
        RECT 87.030 93.520 87.990 93.750 ;
        RECT 88.130 93.595 95.905 94.395 ;
        RECT 96.155 93.750 97.005 95.170 ;
        RECT 88.130 93.320 88.580 93.595 ;
        RECT 86.030 84.295 87.855 93.320 ;
        RECT 88.030 84.295 88.580 93.320 ;
        RECT 89.055 84.295 89.855 93.320 ;
        RECT 90.330 84.295 91.130 93.595 ;
        RECT 91.630 84.295 92.430 93.320 ;
        RECT 92.930 84.295 93.730 93.595 ;
        RECT 95.480 93.320 95.905 93.595 ;
        RECT 96.060 93.520 97.020 93.750 ;
        RECT 97.255 93.320 98.030 95.620 ;
        RECT 94.205 84.295 95.005 93.320 ;
        RECT 95.480 84.295 96.280 93.320 ;
        RECT 97.105 93.315 98.030 93.320 ;
        RECT 97.070 84.315 98.030 93.315 ;
        RECT 97.105 84.295 98.030 84.315 ;
        RECT 99.355 95.620 111.355 95.645 ;
        RECT 99.355 93.320 100.105 95.620 ;
        RECT 100.355 93.750 101.205 95.170 ;
        RECT 101.555 94.820 109.130 95.620 ;
        RECT 100.355 93.520 101.315 93.750 ;
        RECT 101.455 93.595 109.230 94.395 ;
        RECT 109.480 93.750 110.330 95.170 ;
        RECT 101.455 93.320 101.905 93.595 ;
        RECT 99.355 84.295 101.180 93.320 ;
        RECT 101.355 84.295 101.905 93.320 ;
        RECT 102.380 84.295 103.180 93.320 ;
        RECT 103.655 84.295 104.455 93.595 ;
        RECT 104.955 84.295 105.755 93.320 ;
        RECT 106.255 84.295 107.055 93.595 ;
        RECT 108.805 93.320 109.230 93.595 ;
        RECT 109.385 93.520 110.345 93.750 ;
        RECT 110.580 93.320 111.355 95.620 ;
        RECT 107.530 84.295 108.330 93.320 ;
        RECT 108.805 84.295 109.605 93.320 ;
        RECT 110.430 93.315 111.355 93.320 ;
        RECT 110.395 84.315 111.355 93.315 ;
        RECT 110.430 84.295 111.355 84.315 ;
        RECT 112.680 95.595 122.105 95.645 ;
        RECT 112.680 93.320 113.405 95.595 ;
        RECT 113.680 93.750 114.530 95.170 ;
        RECT 114.880 94.670 119.880 95.595 ;
        RECT 113.680 93.520 114.640 93.750 ;
        RECT 114.780 93.595 119.980 94.395 ;
        RECT 120.180 93.750 121.030 95.170 ;
        RECT 114.780 93.320 115.205 93.595 ;
        RECT 112.680 84.295 114.505 93.320 ;
        RECT 114.680 84.295 115.205 93.320 ;
        RECT 115.705 84.295 116.505 93.320 ;
        RECT 116.980 84.295 117.780 93.595 ;
        RECT 119.555 93.320 119.980 93.595 ;
        RECT 120.130 93.520 121.090 93.750 ;
        RECT 121.305 93.320 122.105 95.595 ;
        RECT 118.255 84.295 119.055 93.320 ;
        RECT 119.555 84.295 120.355 93.320 ;
        RECT 121.180 93.315 122.105 93.320 ;
        RECT 121.140 84.315 122.105 93.315 ;
        RECT 121.155 84.295 122.105 84.315 ;
        RECT 123.430 95.620 135.430 95.645 ;
        RECT 123.430 93.320 124.180 95.620 ;
        RECT 124.430 93.750 125.280 95.170 ;
        RECT 125.630 94.820 133.205 95.620 ;
        RECT 124.430 93.520 125.390 93.750 ;
        RECT 125.530 93.595 133.305 94.395 ;
        RECT 133.555 93.750 134.405 95.170 ;
        RECT 125.530 93.320 125.980 93.595 ;
        RECT 123.430 84.295 125.255 93.320 ;
        RECT 125.430 84.295 125.980 93.320 ;
        RECT 126.455 84.295 127.255 93.320 ;
        RECT 127.730 84.295 128.530 93.595 ;
        RECT 129.030 84.295 129.830 93.320 ;
        RECT 130.330 84.295 131.130 93.595 ;
        RECT 132.880 93.320 133.305 93.595 ;
        RECT 133.460 93.520 134.420 93.750 ;
        RECT 134.655 93.320 135.430 95.620 ;
        RECT 131.605 84.295 132.405 93.320 ;
        RECT 132.880 84.295 133.680 93.320 ;
        RECT 134.505 93.315 135.430 93.320 ;
        RECT 134.470 84.315 135.430 93.315 ;
        RECT 134.505 84.295 135.430 84.315 ;
        RECT 136.755 95.620 148.755 95.645 ;
        RECT 136.755 93.320 137.505 95.620 ;
        RECT 137.755 93.750 138.605 95.170 ;
        RECT 138.955 94.820 146.530 95.620 ;
        RECT 137.755 93.520 138.715 93.750 ;
        RECT 138.855 93.595 146.630 94.395 ;
        RECT 146.880 93.750 147.730 95.170 ;
        RECT 138.855 93.320 139.305 93.595 ;
        RECT 136.755 84.295 138.580 93.320 ;
        RECT 138.755 84.295 139.305 93.320 ;
        RECT 139.780 84.295 140.580 93.320 ;
        RECT 141.055 84.295 141.855 93.595 ;
        RECT 142.355 84.295 143.155 93.320 ;
        RECT 143.655 84.295 144.455 93.595 ;
        RECT 146.205 93.320 146.630 93.595 ;
        RECT 146.785 93.520 147.745 93.750 ;
        RECT 147.980 93.320 148.755 95.620 ;
        RECT 144.930 84.295 145.730 93.320 ;
        RECT 146.205 84.295 147.005 93.320 ;
        RECT 147.830 93.315 148.755 93.320 ;
        RECT 147.795 84.315 148.755 93.315 ;
        RECT 147.830 84.295 148.755 84.315 ;
        RECT 150.080 95.620 162.080 95.645 ;
        RECT 150.080 93.320 150.830 95.620 ;
        RECT 151.080 93.750 151.930 95.170 ;
        RECT 152.280 94.820 159.855 95.620 ;
        RECT 151.080 93.520 152.040 93.750 ;
        RECT 152.180 93.595 159.955 94.395 ;
        RECT 160.205 93.750 161.055 95.170 ;
        RECT 152.180 93.320 152.630 93.595 ;
        RECT 150.080 84.295 151.905 93.320 ;
        RECT 152.080 84.295 152.630 93.320 ;
        RECT 153.105 84.295 153.905 93.320 ;
        RECT 154.380 84.295 155.180 93.595 ;
        RECT 155.680 84.295 156.480 93.320 ;
        RECT 156.980 84.295 157.780 93.595 ;
        RECT 159.530 93.320 159.955 93.595 ;
        RECT 160.110 93.520 161.070 93.750 ;
        RECT 161.305 93.320 162.080 95.620 ;
        RECT 158.255 84.295 159.055 93.320 ;
        RECT 159.530 84.295 160.330 93.320 ;
        RECT 161.155 93.315 162.080 93.320 ;
        RECT 161.120 84.315 162.080 93.315 ;
        RECT 161.155 84.295 162.080 84.315 ;
        RECT 163.405 95.620 175.405 95.645 ;
        RECT 163.405 93.320 164.155 95.620 ;
        RECT 164.405 93.750 165.255 95.170 ;
        RECT 165.605 94.820 173.180 95.620 ;
        RECT 164.405 93.520 165.365 93.750 ;
        RECT 165.505 93.595 173.280 94.395 ;
        RECT 173.530 93.750 174.380 95.170 ;
        RECT 165.505 93.320 165.955 93.595 ;
        RECT 163.405 84.295 165.230 93.320 ;
        RECT 165.405 84.295 165.955 93.320 ;
        RECT 166.430 84.295 167.230 93.320 ;
        RECT 167.705 84.295 168.505 93.595 ;
        RECT 169.005 84.295 169.805 93.320 ;
        RECT 170.305 84.295 171.105 93.595 ;
        RECT 172.855 93.320 173.280 93.595 ;
        RECT 173.435 93.520 174.395 93.750 ;
        RECT 174.630 93.320 175.405 95.620 ;
        RECT 171.580 84.295 172.380 93.320 ;
        RECT 172.855 84.295 173.655 93.320 ;
        RECT 174.480 93.315 175.405 93.320 ;
        RECT 174.445 84.315 175.405 93.315 ;
        RECT 174.480 84.295 175.405 84.315 ;
        RECT 176.730 95.620 188.730 95.645 ;
        RECT 176.730 93.320 177.480 95.620 ;
        RECT 177.730 93.750 178.580 95.170 ;
        RECT 178.930 94.820 186.505 95.620 ;
        RECT 177.730 93.520 178.690 93.750 ;
        RECT 178.830 93.595 186.605 94.395 ;
        RECT 186.855 93.750 187.705 95.170 ;
        RECT 178.830 93.320 179.280 93.595 ;
        RECT 176.730 84.295 178.555 93.320 ;
        RECT 178.730 84.295 179.280 93.320 ;
        RECT 179.755 84.295 180.555 93.320 ;
        RECT 181.030 84.295 181.830 93.595 ;
        RECT 182.330 84.295 183.130 93.320 ;
        RECT 183.630 84.295 184.430 93.595 ;
        RECT 186.180 93.320 186.605 93.595 ;
        RECT 186.760 93.520 187.720 93.750 ;
        RECT 187.955 93.320 188.730 95.620 ;
        RECT 184.905 84.295 185.705 93.320 ;
        RECT 186.180 84.295 186.980 93.320 ;
        RECT 187.805 93.315 188.730 93.320 ;
        RECT 187.770 84.315 188.730 93.315 ;
        RECT 187.805 84.295 188.730 84.315 ;
        RECT 190.055 95.595 199.480 95.645 ;
        RECT 190.055 93.320 190.780 95.595 ;
        RECT 191.055 93.750 191.905 95.170 ;
        RECT 192.255 94.670 197.255 95.595 ;
        RECT 191.055 93.520 192.015 93.750 ;
        RECT 192.155 93.595 197.355 94.395 ;
        RECT 197.555 93.750 198.405 95.170 ;
        RECT 192.155 93.320 192.580 93.595 ;
        RECT 190.055 84.295 191.880 93.320 ;
        RECT 192.055 84.295 192.580 93.320 ;
        RECT 193.080 84.295 193.880 93.320 ;
        RECT 194.355 84.295 195.155 93.595 ;
        RECT 196.930 93.320 197.355 93.595 ;
        RECT 197.505 93.520 198.465 93.750 ;
        RECT 198.680 93.320 199.480 95.595 ;
        RECT 195.630 84.295 196.430 93.320 ;
        RECT 196.930 84.295 197.730 93.320 ;
        RECT 198.555 93.315 199.480 93.320 ;
        RECT 198.515 84.315 199.480 93.315 ;
        RECT 198.530 84.295 199.480 84.315 ;
        RECT 200.805 95.620 212.805 95.645 ;
        RECT 200.805 93.320 201.555 95.620 ;
        RECT 201.805 93.750 202.655 95.170 ;
        RECT 203.005 94.820 210.580 95.620 ;
        RECT 201.805 93.520 202.765 93.750 ;
        RECT 202.905 93.595 210.680 94.395 ;
        RECT 210.930 93.750 211.780 95.170 ;
        RECT 202.905 93.320 203.355 93.595 ;
        RECT 200.805 84.295 202.630 93.320 ;
        RECT 202.805 84.295 203.355 93.320 ;
        RECT 203.830 84.295 204.630 93.320 ;
        RECT 205.105 84.295 205.905 93.595 ;
        RECT 206.405 84.295 207.205 93.320 ;
        RECT 207.705 84.295 208.505 93.595 ;
        RECT 210.255 93.320 210.680 93.595 ;
        RECT 210.835 93.520 211.795 93.750 ;
        RECT 212.030 93.320 212.805 95.620 ;
        RECT 208.980 84.295 209.780 93.320 ;
        RECT 210.255 84.295 211.055 93.320 ;
        RECT 211.880 93.315 212.805 93.320 ;
        RECT 211.845 84.315 212.805 93.315 ;
        RECT 211.880 84.295 212.805 84.315 ;
        RECT 214.130 95.620 226.130 95.645 ;
        RECT 214.130 93.320 214.880 95.620 ;
        RECT 215.130 93.750 215.980 95.170 ;
        RECT 216.330 94.820 223.905 95.620 ;
        RECT 215.130 93.520 216.090 93.750 ;
        RECT 216.230 93.595 224.005 94.395 ;
        RECT 224.255 93.750 225.105 95.170 ;
        RECT 216.230 93.320 216.680 93.595 ;
        RECT 214.130 84.295 215.955 93.320 ;
        RECT 216.130 84.295 216.680 93.320 ;
        RECT 217.155 84.295 217.955 93.320 ;
        RECT 218.430 84.295 219.230 93.595 ;
        RECT 219.730 84.295 220.530 93.320 ;
        RECT 221.030 84.295 221.830 93.595 ;
        RECT 223.580 93.320 224.005 93.595 ;
        RECT 224.160 93.520 225.120 93.750 ;
        RECT 225.355 93.320 226.130 95.620 ;
        RECT 222.305 84.295 223.105 93.320 ;
        RECT 223.580 84.295 224.380 93.320 ;
        RECT 225.205 93.315 226.130 93.320 ;
        RECT 225.170 84.315 226.130 93.315 ;
        RECT 225.205 84.295 226.130 84.315 ;
        RECT 226.800 89.700 228.050 97.100 ;
        RECT 228.675 114.075 273.400 114.675 ;
        RECT 228.675 90.150 229.275 114.075 ;
        RECT 275.775 111.700 276.375 169.700 ;
        RECT 230.000 111.100 276.375 111.700 ;
        RECT 230.000 100.475 230.600 111.100 ;
        RECT 240.650 106.350 243.525 106.500 ;
        RECT 231.050 105.495 266.400 106.350 ;
        RECT 231.045 105.150 266.400 105.495 ;
        RECT 231.045 105.145 234.650 105.150 ;
        RECT 235.645 105.145 248.450 105.150 ;
        RECT 231.050 105.125 234.650 105.145 ;
        RECT 231.050 104.400 232.050 105.125 ;
        RECT 233.650 104.945 234.650 105.125 ;
        RECT 233.645 104.620 234.650 104.945 ;
        RECT 233.650 104.400 234.650 104.620 ;
        RECT 231.050 104.395 232.275 104.400 ;
        RECT 231.050 101.400 232.480 104.395 ;
        RECT 232.675 101.400 233.025 104.400 ;
        RECT 233.425 104.395 234.650 104.400 ;
        RECT 233.210 101.400 234.650 104.395 ;
        RECT 235.650 105.125 248.450 105.145 ;
        RECT 235.650 104.400 236.650 105.125 ;
        RECT 238.250 104.945 241.525 105.125 ;
        RECT 242.575 104.945 245.850 105.125 ;
        RECT 247.450 104.945 248.450 105.125 ;
        RECT 238.245 104.625 241.525 104.945 ;
        RECT 238.245 104.620 241.250 104.625 ;
        RECT 242.570 104.620 245.850 104.945 ;
        RECT 247.445 104.620 248.450 104.945 ;
        RECT 238.250 104.400 241.250 104.620 ;
        RECT 242.850 104.400 245.850 104.620 ;
        RECT 247.450 104.400 248.450 104.620 ;
        RECT 235.650 104.395 236.875 104.400 ;
        RECT 235.650 101.400 237.080 104.395 ;
        RECT 237.275 101.400 237.625 104.400 ;
        RECT 238.025 104.395 241.475 104.400 ;
        RECT 237.810 101.400 241.680 104.395 ;
        RECT 241.875 101.400 242.225 104.400 ;
        RECT 242.625 104.395 246.075 104.400 ;
        RECT 242.410 101.400 246.280 104.395 ;
        RECT 246.475 101.400 246.825 104.400 ;
        RECT 247.225 104.395 248.450 104.400 ;
        RECT 247.010 101.400 248.450 104.395 ;
        RECT 249.450 104.950 250.450 105.150 ;
        RECT 249.450 104.625 250.455 104.950 ;
        RECT 249.450 104.400 250.450 104.625 ;
        RECT 249.450 101.400 250.880 104.400 ;
        RECT 251.075 101.400 251.400 104.400 ;
        RECT 251.600 101.400 251.850 105.150 ;
        RECT 252.050 101.400 252.375 104.400 ;
        RECT 252.550 101.400 252.800 105.150 ;
        RECT 253.950 105.000 266.400 105.150 ;
        RECT 253.950 104.400 254.950 105.000 ;
        RECT 253.000 101.400 253.325 104.400 ;
        RECT 253.530 101.400 254.950 104.400 ;
        RECT 231.770 101.395 232.000 101.400 ;
        RECT 232.250 101.395 232.480 101.400 ;
        RECT 232.730 101.395 232.960 101.400 ;
        RECT 233.210 101.395 233.440 101.400 ;
        RECT 233.690 101.395 233.920 101.400 ;
        RECT 236.370 101.395 236.600 101.400 ;
        RECT 236.850 101.395 237.080 101.400 ;
        RECT 237.330 101.395 237.560 101.400 ;
        RECT 237.810 101.395 238.040 101.400 ;
        RECT 238.290 101.395 238.520 101.400 ;
        RECT 240.970 101.395 241.200 101.400 ;
        RECT 241.450 101.395 241.680 101.400 ;
        RECT 241.930 101.395 242.160 101.400 ;
        RECT 242.410 101.395 242.640 101.400 ;
        RECT 242.890 101.395 243.120 101.400 ;
        RECT 245.570 101.395 245.800 101.400 ;
        RECT 246.050 101.395 246.280 101.400 ;
        RECT 246.530 101.395 246.760 101.400 ;
        RECT 247.010 101.395 247.240 101.400 ;
        RECT 247.490 101.395 247.720 101.400 ;
        RECT 232.450 101.195 233.250 101.200 ;
        RECT 237.050 101.195 237.850 101.200 ;
        RECT 242.100 101.195 242.475 101.200 ;
        RECT 246.250 101.195 247.050 101.200 ;
        RECT 232.445 100.820 233.250 101.195 ;
        RECT 237.045 100.820 237.850 101.195 ;
        RECT 242.095 100.820 242.475 101.195 ;
        RECT 246.245 100.820 247.050 101.195 ;
        RECT 232.450 100.475 233.250 100.820 ;
        RECT 237.050 100.475 237.850 100.820 ;
        RECT 242.100 100.475 242.475 100.820 ;
        RECT 246.250 100.475 247.050 100.820 ;
        RECT 250.825 100.825 253.580 101.200 ;
        RECT 250.825 100.475 253.575 100.825 ;
        RECT 230.000 99.875 233.250 100.475 ;
        RECT 234.900 99.875 237.850 100.475 ;
        RECT 239.500 99.875 242.475 100.475 ;
        RECT 244.775 99.875 247.050 100.475 ;
        RECT 248.700 99.875 253.575 100.475 ;
        RECT 230.000 91.175 230.600 99.875 ;
        RECT 232.450 99.200 233.250 99.875 ;
        RECT 237.050 99.200 237.850 99.875 ;
        RECT 242.100 99.200 242.475 99.875 ;
        RECT 246.250 99.200 247.050 99.875 ;
        RECT 250.825 99.525 253.575 99.875 ;
        RECT 250.825 99.200 253.580 99.525 ;
        RECT 256.625 99.450 271.250 99.800 ;
        RECT 231.050 98.000 232.485 99.000 ;
        RECT 232.675 98.000 233.025 99.000 ;
        RECT 233.215 98.000 237.085 99.000 ;
        RECT 237.275 98.000 237.625 99.000 ;
        RECT 237.815 98.000 239.250 99.000 ;
        RECT 231.050 97.300 232.050 98.000 ;
        RECT 233.650 97.300 236.650 98.000 ;
        RECT 238.250 97.300 239.250 98.000 ;
        RECT 240.250 98.000 241.685 99.000 ;
        RECT 241.875 98.000 242.225 99.000 ;
        RECT 242.415 98.000 243.850 99.000 ;
        RECT 240.250 97.800 241.250 98.000 ;
        RECT 242.850 97.800 243.850 98.000 ;
        RECT 240.250 97.300 241.525 97.800 ;
        RECT 242.575 97.300 243.850 97.800 ;
        RECT 244.850 98.000 246.285 99.000 ;
        RECT 246.475 98.000 246.825 99.000 ;
        RECT 247.015 98.000 250.880 99.000 ;
        RECT 251.075 98.000 251.400 99.000 ;
        RECT 244.850 97.300 245.850 98.000 ;
        RECT 247.450 97.975 250.880 98.000 ;
        RECT 247.450 97.300 250.875 97.975 ;
        RECT 251.600 97.300 251.850 99.000 ;
        RECT 252.050 98.000 252.375 99.000 ;
        RECT 252.550 97.300 252.800 99.000 ;
        RECT 253.000 98.000 253.325 99.000 ;
        RECT 253.525 97.300 254.950 99.000 ;
        RECT 256.625 98.900 271.250 99.275 ;
        RECT 231.050 96.950 254.955 97.300 ;
        RECT 231.050 96.200 233.700 96.205 ;
        RECT 231.050 95.850 254.955 96.200 ;
        RECT 231.050 92.100 231.425 95.850 ;
        RECT 231.950 95.300 232.800 95.680 ;
        RECT 231.775 91.175 232.025 95.125 ;
        RECT 232.200 92.100 232.550 95.125 ;
        RECT 232.725 91.175 232.975 95.125 ;
        RECT 233.325 92.100 233.700 95.850 ;
        RECT 235.645 95.845 248.450 95.850 ;
        RECT 235.650 95.825 248.450 95.845 ;
        RECT 235.650 95.100 236.650 95.825 ;
        RECT 238.250 95.645 241.525 95.825 ;
        RECT 242.575 95.645 245.850 95.825 ;
        RECT 247.450 95.645 248.450 95.825 ;
        RECT 238.245 95.325 241.525 95.645 ;
        RECT 238.245 95.320 241.250 95.325 ;
        RECT 242.570 95.320 245.850 95.645 ;
        RECT 247.445 95.320 248.450 95.645 ;
        RECT 238.250 95.100 241.250 95.320 ;
        RECT 242.850 95.100 245.850 95.320 ;
        RECT 247.450 95.100 248.450 95.320 ;
        RECT 235.650 95.095 236.875 95.100 ;
        RECT 235.650 92.100 237.080 95.095 ;
        RECT 237.275 92.100 237.625 95.100 ;
        RECT 238.025 95.095 241.475 95.100 ;
        RECT 237.810 92.100 241.680 95.095 ;
        RECT 241.875 92.100 242.225 95.100 ;
        RECT 242.625 95.095 246.075 95.100 ;
        RECT 242.410 92.100 246.280 95.095 ;
        RECT 246.475 92.100 246.825 95.100 ;
        RECT 247.225 95.095 248.450 95.100 ;
        RECT 247.010 92.100 248.450 95.095 ;
        RECT 249.450 95.650 250.450 95.850 ;
        RECT 249.450 95.325 250.455 95.650 ;
        RECT 249.450 95.100 250.450 95.325 ;
        RECT 249.450 92.100 250.880 95.100 ;
        RECT 251.075 92.100 251.400 95.100 ;
        RECT 251.600 92.100 251.850 95.850 ;
        RECT 252.050 92.100 252.375 95.100 ;
        RECT 252.550 92.100 252.800 95.850 ;
        RECT 253.950 95.100 254.950 95.850 ;
        RECT 253.000 92.100 253.325 95.100 ;
        RECT 253.530 92.100 254.950 95.100 ;
        RECT 256.625 92.100 256.975 98.900 ;
        RECT 257.540 98.895 259.290 98.900 ;
        RECT 268.590 98.895 270.340 98.900 ;
        RECT 257.345 98.625 257.575 98.695 ;
        RECT 257.825 98.625 258.055 98.695 ;
        RECT 258.305 98.625 258.535 98.695 ;
        RECT 258.785 98.625 259.015 98.695 ;
        RECT 259.265 98.625 259.495 98.695 ;
        RECT 259.745 98.625 259.975 98.695 ;
        RECT 257.300 97.450 259.500 98.625 ;
        RECT 259.700 97.450 260.025 98.625 ;
        RECT 257.345 95.695 257.575 97.450 ;
        RECT 257.825 95.695 258.055 97.450 ;
        RECT 258.305 95.695 258.535 97.450 ;
        RECT 258.785 95.695 259.015 97.450 ;
        RECT 259.225 97.425 259.500 97.450 ;
        RECT 259.225 95.700 259.550 97.425 ;
        RECT 259.265 95.695 259.495 95.700 ;
        RECT 259.745 95.695 259.975 97.450 ;
        RECT 260.225 96.875 260.455 98.695 ;
        RECT 260.705 98.625 260.935 98.695 ;
        RECT 260.650 97.450 260.975 98.625 ;
        RECT 260.175 95.700 260.500 96.875 ;
        RECT 260.225 95.695 260.455 95.700 ;
        RECT 260.705 95.695 260.935 97.450 ;
        RECT 261.185 96.875 261.415 98.695 ;
        RECT 261.665 98.625 261.895 98.695 ;
        RECT 261.625 97.450 261.950 98.625 ;
        RECT 261.125 95.700 261.475 96.875 ;
        RECT 261.185 95.695 261.415 95.700 ;
        RECT 261.665 95.695 261.895 97.450 ;
        RECT 262.145 96.875 262.375 98.695 ;
        RECT 262.625 98.625 262.855 98.695 ;
        RECT 262.575 97.450 262.900 98.625 ;
        RECT 262.100 95.700 262.425 96.875 ;
        RECT 262.145 95.695 262.375 95.700 ;
        RECT 262.625 95.695 262.855 97.450 ;
        RECT 263.105 96.875 263.335 98.695 ;
        RECT 263.585 98.625 263.815 98.695 ;
        RECT 263.525 97.450 263.875 98.625 ;
        RECT 263.050 95.700 263.375 96.875 ;
        RECT 263.105 95.695 263.335 95.700 ;
        RECT 263.585 95.695 263.815 97.450 ;
        RECT 264.065 96.875 264.295 98.695 ;
        RECT 264.545 98.625 264.775 98.695 ;
        RECT 264.500 97.450 264.825 98.625 ;
        RECT 264.025 95.700 264.350 96.875 ;
        RECT 264.065 95.695 264.295 95.700 ;
        RECT 264.545 95.695 264.775 97.450 ;
        RECT 265.025 96.875 265.255 98.695 ;
        RECT 265.505 98.625 265.735 98.695 ;
        RECT 265.450 97.450 265.775 98.625 ;
        RECT 264.975 95.700 265.300 96.875 ;
        RECT 265.025 95.695 265.255 95.700 ;
        RECT 265.505 95.695 265.735 97.450 ;
        RECT 265.985 96.875 266.215 98.695 ;
        RECT 266.465 98.625 266.695 98.695 ;
        RECT 266.425 97.450 266.750 98.625 ;
        RECT 265.925 95.700 266.250 96.875 ;
        RECT 265.985 95.695 266.215 95.700 ;
        RECT 266.465 95.695 266.695 97.450 ;
        RECT 266.945 96.875 267.175 98.695 ;
        RECT 267.425 98.625 267.655 98.695 ;
        RECT 267.375 97.450 267.700 98.625 ;
        RECT 266.900 95.700 267.225 96.875 ;
        RECT 266.945 95.695 267.175 95.700 ;
        RECT 267.425 95.695 267.655 97.450 ;
        RECT 267.905 96.875 268.135 98.695 ;
        RECT 268.385 98.625 268.615 98.695 ;
        RECT 268.865 98.625 269.095 98.695 ;
        RECT 269.345 98.625 269.575 98.695 ;
        RECT 269.825 98.625 270.055 98.695 ;
        RECT 270.305 98.625 270.535 98.695 ;
        RECT 268.325 97.450 270.575 98.625 ;
        RECT 267.850 95.700 268.175 96.875 ;
        RECT 267.905 95.695 268.135 95.700 ;
        RECT 268.385 95.695 268.615 97.450 ;
        RECT 268.865 95.695 269.095 97.450 ;
        RECT 269.345 95.695 269.575 97.450 ;
        RECT 269.825 95.695 270.055 97.450 ;
        RECT 270.305 95.695 270.535 97.450 ;
        RECT 257.525 93.500 270.350 95.500 ;
        RECT 257.345 92.650 257.575 93.300 ;
        RECT 257.825 92.650 258.055 93.300 ;
        RECT 258.305 92.650 258.535 93.300 ;
        RECT 258.785 92.650 259.015 93.300 ;
        RECT 259.225 92.675 259.550 93.300 ;
        RECT 259.225 92.650 259.525 92.675 ;
        RECT 259.745 92.650 259.975 93.300 ;
        RECT 260.175 92.900 260.500 93.300 ;
        RECT 257.300 92.250 259.525 92.650 ;
        RECT 259.700 92.250 260.025 92.650 ;
        RECT 260.225 92.300 260.455 92.900 ;
        RECT 260.705 92.650 260.935 93.300 ;
        RECT 261.125 92.900 261.475 93.300 ;
        RECT 260.650 92.250 261.000 92.650 ;
        RECT 261.185 92.300 261.415 92.900 ;
        RECT 261.665 92.650 261.895 93.300 ;
        RECT 262.100 92.900 262.425 93.300 ;
        RECT 261.625 92.250 261.950 92.650 ;
        RECT 262.145 92.300 262.375 92.900 ;
        RECT 262.625 92.650 262.855 93.300 ;
        RECT 263.050 92.900 263.375 93.300 ;
        RECT 262.575 92.250 262.900 92.650 ;
        RECT 263.105 92.300 263.335 92.900 ;
        RECT 263.585 92.650 263.815 93.300 ;
        RECT 264.025 92.900 264.350 93.300 ;
        RECT 263.525 92.250 263.875 92.650 ;
        RECT 264.065 92.300 264.295 92.900 ;
        RECT 264.545 92.650 264.775 93.300 ;
        RECT 264.975 92.900 265.300 93.300 ;
        RECT 264.500 92.250 264.825 92.650 ;
        RECT 265.025 92.300 265.255 92.900 ;
        RECT 265.505 92.650 265.735 93.300 ;
        RECT 265.925 92.900 266.275 93.300 ;
        RECT 265.450 92.250 265.800 92.650 ;
        RECT 265.985 92.300 266.215 92.900 ;
        RECT 266.465 92.650 266.695 93.300 ;
        RECT 266.900 92.900 267.225 93.300 ;
        RECT 266.425 92.250 266.750 92.650 ;
        RECT 266.945 92.300 267.175 92.900 ;
        RECT 267.425 92.650 267.655 93.300 ;
        RECT 267.850 92.900 268.200 93.300 ;
        RECT 267.375 92.250 267.700 92.650 ;
        RECT 267.905 92.300 268.135 92.900 ;
        RECT 268.385 92.650 268.615 93.300 ;
        RECT 268.865 92.650 269.095 93.300 ;
        RECT 269.345 92.650 269.575 93.300 ;
        RECT 269.825 92.650 270.055 93.300 ;
        RECT 270.305 92.650 270.535 93.300 ;
        RECT 268.325 92.250 270.575 92.650 ;
        RECT 270.900 92.100 271.250 98.900 ;
        RECT 236.370 92.095 236.600 92.100 ;
        RECT 236.850 92.095 237.080 92.100 ;
        RECT 237.330 92.095 237.560 92.100 ;
        RECT 237.810 92.095 238.040 92.100 ;
        RECT 238.290 92.095 238.520 92.100 ;
        RECT 240.970 92.095 241.200 92.100 ;
        RECT 241.450 92.095 241.680 92.100 ;
        RECT 241.930 92.095 242.160 92.100 ;
        RECT 242.410 92.095 242.640 92.100 ;
        RECT 242.890 92.095 243.120 92.100 ;
        RECT 245.570 92.095 245.800 92.100 ;
        RECT 246.050 92.095 246.280 92.100 ;
        RECT 246.530 92.095 246.760 92.100 ;
        RECT 247.010 92.095 247.240 92.100 ;
        RECT 247.490 92.095 247.720 92.100 ;
        RECT 237.050 91.895 237.850 91.900 ;
        RECT 242.100 91.895 242.475 91.900 ;
        RECT 246.250 91.895 247.050 91.900 ;
        RECT 230.000 90.575 232.975 91.175 ;
        RECT 226.800 88.000 231.425 89.700 ;
        RECT 231.775 88.700 232.025 90.575 ;
        RECT 232.200 88.700 232.550 89.700 ;
        RECT 232.725 88.700 232.975 90.575 ;
        RECT 233.325 89.700 233.700 91.850 ;
        RECT 237.045 91.520 237.850 91.895 ;
        RECT 242.095 91.520 242.475 91.895 ;
        RECT 246.245 91.520 247.050 91.895 ;
        RECT 237.050 91.175 237.850 91.520 ;
        RECT 242.100 91.175 242.475 91.520 ;
        RECT 246.250 91.175 247.050 91.520 ;
        RECT 250.825 91.525 253.580 91.900 ;
        RECT 256.625 91.775 271.250 92.100 ;
        RECT 250.825 91.175 253.575 91.525 ;
        RECT 256.625 91.250 271.250 91.600 ;
        RECT 234.900 90.575 237.850 91.175 ;
        RECT 239.500 90.575 242.475 91.175 ;
        RECT 244.775 90.575 247.050 91.175 ;
        RECT 248.700 90.575 253.575 91.175 ;
        RECT 237.050 89.900 237.850 90.575 ;
        RECT 242.100 89.900 242.475 90.575 ;
        RECT 246.250 89.900 247.050 90.575 ;
        RECT 250.825 90.225 253.575 90.575 ;
        RECT 250.825 89.900 253.580 90.225 ;
        RECT 233.325 88.700 237.085 89.700 ;
        RECT 237.275 88.700 237.625 89.700 ;
        RECT 237.815 88.700 239.250 89.700 ;
        RECT 231.950 88.175 232.800 88.500 ;
        RECT 233.325 88.000 236.650 88.700 ;
        RECT 238.250 88.000 239.250 88.700 ;
        RECT 240.250 88.700 241.685 89.700 ;
        RECT 241.875 88.700 242.225 89.700 ;
        RECT 242.415 88.700 243.850 89.700 ;
        RECT 240.250 88.500 241.250 88.700 ;
        RECT 242.850 88.500 243.850 88.700 ;
        RECT 240.250 88.000 241.525 88.500 ;
        RECT 242.575 88.000 243.850 88.500 ;
        RECT 244.850 88.700 246.285 89.700 ;
        RECT 246.475 88.700 246.825 89.700 ;
        RECT 247.015 88.700 250.880 89.700 ;
        RECT 251.075 88.700 251.400 89.700 ;
        RECT 244.850 88.000 245.850 88.700 ;
        RECT 247.450 88.675 250.880 88.700 ;
        RECT 247.450 88.000 250.875 88.675 ;
        RECT 251.600 88.000 251.850 89.700 ;
        RECT 252.050 88.700 252.375 89.700 ;
        RECT 252.550 88.000 252.800 89.700 ;
        RECT 253.000 88.700 253.325 89.700 ;
        RECT 253.525 88.150 254.950 89.700 ;
        RECT 253.525 88.000 261.450 88.150 ;
        RECT 226.800 86.800 261.450 88.000 ;
        RECT 77.570 84.070 78.530 84.110 ;
        RECT 78.860 84.070 79.820 84.110 ;
        RECT 80.150 84.070 81.110 84.110 ;
        RECT 81.440 84.070 82.400 84.110 ;
        RECT 88.320 84.070 89.280 84.110 ;
        RECT 89.610 84.095 90.570 84.110 ;
        RECT 90.900 84.095 91.860 84.110 ;
        RECT 89.610 84.070 91.860 84.095 ;
        RECT 92.190 84.070 93.150 84.110 ;
        RECT 93.480 84.070 94.440 84.110 ;
        RECT 94.770 84.070 95.730 84.110 ;
        RECT 77.570 83.895 82.430 84.070 ;
        RECT 88.320 83.895 95.730 84.070 ;
        RECT 101.645 84.070 102.605 84.110 ;
        RECT 102.935 84.095 103.895 84.110 ;
        RECT 104.225 84.095 105.185 84.110 ;
        RECT 102.935 84.070 105.185 84.095 ;
        RECT 105.515 84.070 106.475 84.110 ;
        RECT 106.805 84.070 107.765 84.110 ;
        RECT 108.095 84.070 109.055 84.110 ;
        RECT 101.645 83.895 109.055 84.070 ;
        RECT 114.970 84.070 115.930 84.110 ;
        RECT 116.260 84.070 117.220 84.110 ;
        RECT 117.550 84.070 118.510 84.110 ;
        RECT 118.840 84.070 119.800 84.110 ;
        RECT 125.720 84.070 126.680 84.110 ;
        RECT 127.010 84.095 127.970 84.110 ;
        RECT 128.300 84.095 129.260 84.110 ;
        RECT 127.010 84.070 129.260 84.095 ;
        RECT 129.590 84.070 130.550 84.110 ;
        RECT 130.880 84.070 131.840 84.110 ;
        RECT 132.170 84.070 133.130 84.110 ;
        RECT 114.970 84.045 119.830 84.070 ;
        RECT 114.970 83.895 120.805 84.045 ;
        RECT 125.720 83.895 133.130 84.070 ;
        RECT 139.045 84.070 140.005 84.110 ;
        RECT 140.335 84.095 141.295 84.110 ;
        RECT 141.625 84.095 142.585 84.110 ;
        RECT 140.335 84.070 142.585 84.095 ;
        RECT 142.915 84.070 143.875 84.110 ;
        RECT 144.205 84.070 145.165 84.110 ;
        RECT 145.495 84.070 146.455 84.110 ;
        RECT 139.045 83.895 146.455 84.070 ;
        RECT 152.370 84.070 153.330 84.110 ;
        RECT 153.660 84.095 154.620 84.110 ;
        RECT 154.950 84.095 155.910 84.110 ;
        RECT 153.660 84.070 155.910 84.095 ;
        RECT 156.240 84.070 157.200 84.110 ;
        RECT 157.530 84.070 158.490 84.110 ;
        RECT 158.820 84.070 159.780 84.110 ;
        RECT 152.370 83.895 159.780 84.070 ;
        RECT 165.695 84.070 166.655 84.110 ;
        RECT 166.985 84.095 167.945 84.110 ;
        RECT 168.275 84.095 169.235 84.110 ;
        RECT 166.985 84.070 169.235 84.095 ;
        RECT 169.565 84.070 170.525 84.110 ;
        RECT 170.855 84.070 171.815 84.110 ;
        RECT 172.145 84.070 173.105 84.110 ;
        RECT 165.695 83.895 173.105 84.070 ;
        RECT 179.020 84.070 179.980 84.110 ;
        RECT 180.310 84.095 181.270 84.110 ;
        RECT 181.600 84.095 182.560 84.110 ;
        RECT 180.310 84.070 182.560 84.095 ;
        RECT 182.890 84.070 183.850 84.110 ;
        RECT 184.180 84.070 185.140 84.110 ;
        RECT 185.470 84.070 186.430 84.110 ;
        RECT 179.020 83.895 186.430 84.070 ;
        RECT 192.345 84.070 193.305 84.110 ;
        RECT 193.635 84.070 194.595 84.110 ;
        RECT 194.925 84.070 195.885 84.110 ;
        RECT 196.215 84.070 197.175 84.110 ;
        RECT 203.095 84.070 204.055 84.110 ;
        RECT 204.385 84.095 205.345 84.110 ;
        RECT 205.675 84.095 206.635 84.110 ;
        RECT 204.385 84.070 206.635 84.095 ;
        RECT 206.965 84.070 207.925 84.110 ;
        RECT 208.255 84.070 209.215 84.110 ;
        RECT 209.545 84.070 210.505 84.110 ;
        RECT 192.345 83.895 198.180 84.070 ;
        RECT 203.095 83.895 210.505 84.070 ;
        RECT 216.420 84.070 217.380 84.110 ;
        RECT 217.710 84.095 218.670 84.110 ;
        RECT 219.000 84.095 219.960 84.110 ;
        RECT 217.710 84.070 219.960 84.095 ;
        RECT 220.290 84.070 221.250 84.110 ;
        RECT 221.580 84.070 222.540 84.110 ;
        RECT 222.870 84.070 223.830 84.110 ;
        RECT 216.420 83.895 223.830 84.070 ;
        RECT 72.650 83.745 75.200 83.750 ;
        RECT 77.555 83.745 82.430 83.895 ;
        RECT 72.650 82.500 82.430 83.745 ;
        RECT 75.105 82.495 82.430 82.500 ;
        RECT 77.555 82.345 82.430 82.495 ;
        RECT 85.680 82.345 95.730 83.895 ;
        RECT 99.005 82.345 109.055 83.895 ;
        RECT 110.755 82.345 120.805 83.895 ;
        RECT 123.080 82.345 133.130 83.895 ;
        RECT 136.405 82.345 146.455 83.895 ;
        RECT 149.730 82.345 159.780 83.895 ;
        RECT 163.055 82.345 173.105 83.895 ;
        RECT 176.380 82.345 186.430 83.895 ;
        RECT 189.705 82.345 198.180 83.895 ;
        RECT 200.455 82.345 210.505 83.895 ;
        RECT 213.780 82.345 223.830 83.895 ;
        RECT 77.570 82.170 82.430 82.345 ;
        RECT 88.320 82.170 95.730 82.345 ;
        RECT 77.570 82.130 78.530 82.170 ;
        RECT 78.860 82.130 79.820 82.170 ;
        RECT 80.150 82.130 81.110 82.170 ;
        RECT 81.440 82.130 82.400 82.170 ;
        RECT 88.320 82.130 89.280 82.170 ;
        RECT 89.610 82.145 91.860 82.170 ;
        RECT 89.610 82.130 90.570 82.145 ;
        RECT 90.900 82.130 91.860 82.145 ;
        RECT 92.190 82.130 93.150 82.170 ;
        RECT 93.480 82.130 94.440 82.170 ;
        RECT 94.770 82.130 95.730 82.170 ;
        RECT 101.645 82.170 109.055 82.345 ;
        RECT 101.645 82.130 102.605 82.170 ;
        RECT 102.935 82.145 105.185 82.170 ;
        RECT 102.935 82.130 103.895 82.145 ;
        RECT 104.225 82.130 105.185 82.145 ;
        RECT 105.515 82.130 106.475 82.170 ;
        RECT 106.805 82.130 107.765 82.170 ;
        RECT 108.095 82.130 109.055 82.170 ;
        RECT 114.970 82.170 120.805 82.345 ;
        RECT 125.720 82.170 133.130 82.345 ;
        RECT 114.970 82.130 115.930 82.170 ;
        RECT 116.260 82.130 117.220 82.170 ;
        RECT 117.550 82.130 118.510 82.170 ;
        RECT 118.840 82.130 119.800 82.170 ;
        RECT 125.720 82.130 126.680 82.170 ;
        RECT 127.010 82.145 129.260 82.170 ;
        RECT 127.010 82.130 127.970 82.145 ;
        RECT 128.300 82.130 129.260 82.145 ;
        RECT 129.590 82.130 130.550 82.170 ;
        RECT 130.880 82.130 131.840 82.170 ;
        RECT 132.170 82.130 133.130 82.170 ;
        RECT 139.045 82.170 146.455 82.345 ;
        RECT 139.045 82.130 140.005 82.170 ;
        RECT 140.335 82.145 142.585 82.170 ;
        RECT 140.335 82.130 141.295 82.145 ;
        RECT 141.625 82.130 142.585 82.145 ;
        RECT 142.915 82.130 143.875 82.170 ;
        RECT 144.205 82.130 145.165 82.170 ;
        RECT 145.495 82.130 146.455 82.170 ;
        RECT 152.370 82.170 159.780 82.345 ;
        RECT 152.370 82.130 153.330 82.170 ;
        RECT 153.660 82.145 155.910 82.170 ;
        RECT 153.660 82.130 154.620 82.145 ;
        RECT 154.950 82.130 155.910 82.145 ;
        RECT 156.240 82.130 157.200 82.170 ;
        RECT 157.530 82.130 158.490 82.170 ;
        RECT 158.820 82.130 159.780 82.170 ;
        RECT 165.695 82.170 173.105 82.345 ;
        RECT 165.695 82.130 166.655 82.170 ;
        RECT 166.985 82.145 169.235 82.170 ;
        RECT 166.985 82.130 167.945 82.145 ;
        RECT 168.275 82.130 169.235 82.145 ;
        RECT 169.565 82.130 170.525 82.170 ;
        RECT 170.855 82.130 171.815 82.170 ;
        RECT 172.145 82.130 173.105 82.170 ;
        RECT 179.020 82.170 186.430 82.345 ;
        RECT 179.020 82.130 179.980 82.170 ;
        RECT 180.310 82.145 182.560 82.170 ;
        RECT 180.310 82.130 181.270 82.145 ;
        RECT 181.600 82.130 182.560 82.145 ;
        RECT 182.890 82.130 183.850 82.170 ;
        RECT 184.180 82.130 185.140 82.170 ;
        RECT 185.470 82.130 186.430 82.170 ;
        RECT 192.345 82.170 198.180 82.345 ;
        RECT 203.095 82.170 210.505 82.345 ;
        RECT 192.345 82.130 193.305 82.170 ;
        RECT 193.635 82.130 194.595 82.170 ;
        RECT 194.925 82.130 195.885 82.170 ;
        RECT 196.215 82.130 197.175 82.170 ;
        RECT 203.095 82.130 204.055 82.170 ;
        RECT 204.385 82.145 206.635 82.170 ;
        RECT 204.385 82.130 205.345 82.145 ;
        RECT 205.675 82.130 206.635 82.145 ;
        RECT 206.965 82.130 207.925 82.170 ;
        RECT 208.255 82.130 209.215 82.170 ;
        RECT 209.545 82.130 210.505 82.170 ;
        RECT 216.420 82.170 223.830 82.345 ;
        RECT 216.420 82.130 217.380 82.170 ;
        RECT 217.710 82.145 219.960 82.170 ;
        RECT 217.710 82.130 218.670 82.145 ;
        RECT 219.000 82.130 219.960 82.145 ;
        RECT 220.290 82.130 221.250 82.170 ;
        RECT 221.580 82.130 222.540 82.170 ;
        RECT 222.870 82.130 223.830 82.170 ;
        RECT 226.800 82.000 228.050 86.800 ;
        RECT 226.125 81.995 228.050 82.000 ;
        RECT 75.280 81.925 77.830 81.970 ;
        RECT 75.275 79.025 77.830 81.925 ;
        RECT 75.280 78.695 77.830 79.025 ;
        RECT 78.305 78.970 79.105 81.970 ;
        RECT 79.580 78.695 80.380 81.970 ;
        RECT 80.855 78.970 81.655 81.970 ;
        RECT 82.130 78.695 84.705 81.970 ;
        RECT 75.280 77.625 84.705 78.695 ;
        RECT 75.025 76.695 84.705 77.625 ;
        RECT 86.030 78.970 86.980 81.995 ;
        RECT 97.105 81.970 98.030 81.995 ;
        RECT 87.755 78.970 88.555 81.970 ;
        RECT 89.055 78.970 89.855 81.970 ;
        RECT 86.030 78.945 86.955 78.970 ;
        RECT 86.030 76.720 86.780 78.945 ;
        RECT 87.030 78.580 87.990 78.810 ;
        RECT 88.130 78.695 88.555 78.970 ;
        RECT 90.330 78.695 91.130 81.970 ;
        RECT 91.630 78.970 92.430 81.970 ;
        RECT 92.905 78.695 93.705 81.970 ;
        RECT 94.205 78.970 95.005 81.970 ;
        RECT 95.480 78.970 96.280 81.970 ;
        RECT 97.070 78.970 98.030 81.970 ;
        RECT 95.480 78.695 95.905 78.970 ;
        RECT 87.030 77.170 87.880 78.580 ;
        RECT 88.130 77.895 95.905 78.695 ;
        RECT 96.060 78.580 97.020 78.810 ;
        RECT 88.230 76.720 95.805 77.520 ;
        RECT 96.155 77.170 97.005 78.580 ;
        RECT 97.255 76.720 98.030 78.970 ;
        RECT 86.030 76.695 98.030 76.720 ;
        RECT 99.355 78.970 100.305 81.995 ;
        RECT 110.430 81.970 111.355 81.995 ;
        RECT 101.080 78.970 101.880 81.970 ;
        RECT 102.380 78.970 103.180 81.970 ;
        RECT 99.355 78.945 100.280 78.970 ;
        RECT 99.355 76.720 100.105 78.945 ;
        RECT 100.355 78.580 101.315 78.810 ;
        RECT 101.455 78.695 101.880 78.970 ;
        RECT 103.655 78.695 104.455 81.970 ;
        RECT 104.955 78.970 105.755 81.970 ;
        RECT 106.230 78.695 107.030 81.970 ;
        RECT 107.530 78.970 108.330 81.970 ;
        RECT 108.805 78.970 109.605 81.970 ;
        RECT 110.395 78.970 111.355 81.970 ;
        RECT 108.805 78.695 109.230 78.970 ;
        RECT 100.355 77.170 101.205 78.580 ;
        RECT 101.455 77.895 109.230 78.695 ;
        RECT 109.385 78.580 110.345 78.810 ;
        RECT 101.555 76.720 109.130 77.520 ;
        RECT 109.480 77.170 110.330 78.580 ;
        RECT 110.580 76.720 111.355 78.970 ;
        RECT 99.355 76.695 111.355 76.720 ;
        RECT 112.680 78.945 113.630 81.970 ;
        RECT 114.405 78.970 115.205 81.970 ;
        RECT 115.705 78.970 116.505 81.970 ;
        RECT 112.680 76.695 113.405 78.945 ;
        RECT 113.680 78.580 114.640 78.810 ;
        RECT 114.780 78.695 115.205 78.970 ;
        RECT 116.980 78.695 117.780 81.970 ;
        RECT 118.255 78.970 119.055 81.970 ;
        RECT 119.555 78.970 120.355 81.970 ;
        RECT 121.140 78.970 122.105 81.970 ;
        RECT 119.555 78.695 119.980 78.970 ;
        RECT 121.155 78.945 122.105 78.970 ;
        RECT 113.680 77.170 114.530 78.580 ;
        RECT 114.780 77.895 119.980 78.695 ;
        RECT 120.130 78.580 121.090 78.810 ;
        RECT 114.880 76.695 119.880 77.620 ;
        RECT 120.180 77.170 121.030 78.580 ;
        RECT 121.305 76.695 122.105 78.945 ;
        RECT 123.430 78.970 124.380 81.995 ;
        RECT 134.505 81.970 135.430 81.995 ;
        RECT 125.155 78.970 125.955 81.970 ;
        RECT 126.455 78.970 127.255 81.970 ;
        RECT 123.430 78.945 124.355 78.970 ;
        RECT 123.430 76.720 124.180 78.945 ;
        RECT 124.430 78.580 125.390 78.810 ;
        RECT 125.530 78.695 125.955 78.970 ;
        RECT 127.730 78.695 128.530 81.970 ;
        RECT 129.030 78.970 129.830 81.970 ;
        RECT 130.305 78.695 131.105 81.970 ;
        RECT 131.605 78.970 132.405 81.970 ;
        RECT 132.880 78.970 133.680 81.970 ;
        RECT 134.470 78.970 135.430 81.970 ;
        RECT 132.880 78.695 133.305 78.970 ;
        RECT 124.430 77.170 125.280 78.580 ;
        RECT 125.530 77.895 133.305 78.695 ;
        RECT 133.460 78.580 134.420 78.810 ;
        RECT 125.630 76.720 133.205 77.520 ;
        RECT 133.555 77.170 134.405 78.580 ;
        RECT 134.655 76.720 135.430 78.970 ;
        RECT 123.430 76.695 135.430 76.720 ;
        RECT 136.755 78.970 137.705 81.995 ;
        RECT 147.830 81.970 148.755 81.995 ;
        RECT 138.480 78.970 139.280 81.970 ;
        RECT 139.780 78.970 140.580 81.970 ;
        RECT 136.755 78.945 137.680 78.970 ;
        RECT 136.755 76.720 137.505 78.945 ;
        RECT 137.755 78.580 138.715 78.810 ;
        RECT 138.855 78.695 139.280 78.970 ;
        RECT 141.055 78.695 141.855 81.970 ;
        RECT 142.355 78.970 143.155 81.970 ;
        RECT 143.630 78.695 144.430 81.970 ;
        RECT 144.930 78.970 145.730 81.970 ;
        RECT 146.205 78.970 147.005 81.970 ;
        RECT 147.795 78.970 148.755 81.970 ;
        RECT 146.205 78.695 146.630 78.970 ;
        RECT 137.755 77.170 138.605 78.580 ;
        RECT 138.855 77.895 146.630 78.695 ;
        RECT 146.785 78.580 147.745 78.810 ;
        RECT 138.955 76.720 146.530 77.520 ;
        RECT 146.880 77.170 147.730 78.580 ;
        RECT 147.980 76.720 148.755 78.970 ;
        RECT 136.755 76.695 148.755 76.720 ;
        RECT 150.080 78.970 151.030 81.995 ;
        RECT 161.155 81.970 162.080 81.995 ;
        RECT 151.805 78.970 152.605 81.970 ;
        RECT 153.105 78.970 153.905 81.970 ;
        RECT 150.080 78.945 151.005 78.970 ;
        RECT 150.080 76.720 150.830 78.945 ;
        RECT 151.080 78.580 152.040 78.810 ;
        RECT 152.180 78.695 152.605 78.970 ;
        RECT 154.380 78.695 155.180 81.970 ;
        RECT 155.680 78.970 156.480 81.970 ;
        RECT 156.955 78.695 157.755 81.970 ;
        RECT 158.255 78.970 159.055 81.970 ;
        RECT 159.530 78.970 160.330 81.970 ;
        RECT 161.120 78.970 162.080 81.970 ;
        RECT 159.530 78.695 159.955 78.970 ;
        RECT 151.080 77.170 151.930 78.580 ;
        RECT 152.180 77.895 159.955 78.695 ;
        RECT 160.110 78.580 161.070 78.810 ;
        RECT 152.280 76.720 159.855 77.520 ;
        RECT 160.205 77.170 161.055 78.580 ;
        RECT 161.305 76.720 162.080 78.970 ;
        RECT 150.080 76.695 162.080 76.720 ;
        RECT 163.405 78.970 164.355 81.995 ;
        RECT 174.480 81.970 175.405 81.995 ;
        RECT 165.130 78.970 165.930 81.970 ;
        RECT 166.430 78.970 167.230 81.970 ;
        RECT 163.405 78.945 164.330 78.970 ;
        RECT 163.405 76.720 164.155 78.945 ;
        RECT 164.405 78.580 165.365 78.810 ;
        RECT 165.505 78.695 165.930 78.970 ;
        RECT 167.705 78.695 168.505 81.970 ;
        RECT 169.005 78.970 169.805 81.970 ;
        RECT 170.280 78.695 171.080 81.970 ;
        RECT 171.580 78.970 172.380 81.970 ;
        RECT 172.855 78.970 173.655 81.970 ;
        RECT 174.445 78.970 175.405 81.970 ;
        RECT 172.855 78.695 173.280 78.970 ;
        RECT 164.405 77.170 165.255 78.580 ;
        RECT 165.505 77.895 173.280 78.695 ;
        RECT 173.435 78.580 174.395 78.810 ;
        RECT 165.605 76.720 173.180 77.520 ;
        RECT 173.530 77.170 174.380 78.580 ;
        RECT 174.630 76.720 175.405 78.970 ;
        RECT 163.405 76.695 175.405 76.720 ;
        RECT 176.730 78.970 177.680 81.995 ;
        RECT 187.805 81.970 188.730 81.995 ;
        RECT 178.455 78.970 179.255 81.970 ;
        RECT 179.755 78.970 180.555 81.970 ;
        RECT 176.730 78.945 177.655 78.970 ;
        RECT 176.730 76.720 177.480 78.945 ;
        RECT 177.730 78.580 178.690 78.810 ;
        RECT 178.830 78.695 179.255 78.970 ;
        RECT 181.030 78.695 181.830 81.970 ;
        RECT 182.330 78.970 183.130 81.970 ;
        RECT 183.605 78.695 184.405 81.970 ;
        RECT 184.905 78.970 185.705 81.970 ;
        RECT 186.180 78.970 186.980 81.970 ;
        RECT 187.770 78.970 188.730 81.970 ;
        RECT 186.180 78.695 186.605 78.970 ;
        RECT 177.730 77.170 178.580 78.580 ;
        RECT 178.830 77.895 186.605 78.695 ;
        RECT 186.760 78.580 187.720 78.810 ;
        RECT 178.930 76.720 186.505 77.520 ;
        RECT 186.855 77.170 187.705 78.580 ;
        RECT 187.955 76.720 188.730 78.970 ;
        RECT 176.730 76.695 188.730 76.720 ;
        RECT 190.055 78.945 191.005 81.970 ;
        RECT 191.780 78.970 192.580 81.970 ;
        RECT 193.080 78.970 193.880 81.970 ;
        RECT 190.055 76.695 190.780 78.945 ;
        RECT 191.055 78.580 192.015 78.810 ;
        RECT 192.155 78.695 192.580 78.970 ;
        RECT 194.355 78.695 195.155 81.970 ;
        RECT 195.630 78.970 196.430 81.970 ;
        RECT 196.930 78.970 197.730 81.970 ;
        RECT 198.515 78.970 199.480 81.970 ;
        RECT 196.930 78.695 197.355 78.970 ;
        RECT 198.530 78.945 199.480 78.970 ;
        RECT 191.055 77.170 191.905 78.580 ;
        RECT 192.155 77.895 197.355 78.695 ;
        RECT 197.505 78.580 198.465 78.810 ;
        RECT 192.255 76.695 197.255 77.620 ;
        RECT 197.555 77.170 198.405 78.580 ;
        RECT 198.680 76.695 199.480 78.945 ;
        RECT 200.805 78.970 201.755 81.995 ;
        RECT 211.880 81.970 212.805 81.995 ;
        RECT 202.530 78.970 203.330 81.970 ;
        RECT 203.830 78.970 204.630 81.970 ;
        RECT 200.805 78.945 201.730 78.970 ;
        RECT 200.805 76.720 201.555 78.945 ;
        RECT 201.805 78.580 202.765 78.810 ;
        RECT 202.905 78.695 203.330 78.970 ;
        RECT 205.105 78.695 205.905 81.970 ;
        RECT 206.405 78.970 207.205 81.970 ;
        RECT 207.680 78.695 208.480 81.970 ;
        RECT 208.980 78.970 209.780 81.970 ;
        RECT 210.255 78.970 211.055 81.970 ;
        RECT 211.845 78.970 212.805 81.970 ;
        RECT 210.255 78.695 210.680 78.970 ;
        RECT 201.805 77.170 202.655 78.580 ;
        RECT 202.905 77.895 210.680 78.695 ;
        RECT 210.835 78.580 211.795 78.810 ;
        RECT 203.005 76.720 210.580 77.520 ;
        RECT 210.930 77.170 211.780 78.580 ;
        RECT 212.030 76.720 212.805 78.970 ;
        RECT 200.805 76.695 212.805 76.720 ;
        RECT 214.130 78.970 215.080 81.995 ;
        RECT 225.205 81.970 228.050 81.995 ;
        RECT 215.855 78.970 216.655 81.970 ;
        RECT 217.155 78.970 217.955 81.970 ;
        RECT 214.130 78.945 215.055 78.970 ;
        RECT 214.130 76.720 214.880 78.945 ;
        RECT 215.130 78.580 216.090 78.810 ;
        RECT 216.230 78.695 216.655 78.970 ;
        RECT 218.430 78.695 219.230 81.970 ;
        RECT 219.730 78.970 220.530 81.970 ;
        RECT 221.005 78.695 221.805 81.970 ;
        RECT 222.305 78.970 223.105 81.970 ;
        RECT 223.580 78.970 224.380 81.970 ;
        RECT 225.170 78.970 228.050 81.970 ;
        RECT 223.580 78.695 224.005 78.970 ;
        RECT 215.130 77.170 215.980 78.580 ;
        RECT 216.230 77.895 224.005 78.695 ;
        RECT 224.160 78.580 225.120 78.810 ;
        RECT 216.330 76.720 223.905 77.520 ;
        RECT 224.255 77.170 225.105 78.580 ;
        RECT 225.355 76.720 228.050 78.970 ;
        RECT 214.130 76.695 228.050 76.720 ;
        RECT 75.025 75.950 228.050 76.695 ;
        RECT 75.030 75.945 228.050 75.950 ;
        RECT 111.950 74.635 113.050 74.750 ;
        RECT 97.830 74.600 98.080 74.635 ;
        RECT 98.660 74.600 98.910 74.635 ;
        RECT 99.490 74.600 99.740 74.635 ;
        RECT 100.320 74.600 100.570 74.635 ;
        RECT 101.150 74.600 101.400 74.635 ;
        RECT 101.980 74.600 102.230 74.635 ;
        RECT 102.810 74.600 103.060 74.635 ;
        RECT 103.640 74.600 103.890 74.635 ;
        RECT 104.470 74.600 104.720 74.635 ;
        RECT 105.300 74.600 105.550 74.635 ;
        RECT 106.130 74.600 106.380 74.635 ;
        RECT 106.960 74.600 107.210 74.635 ;
        RECT 107.790 74.600 108.040 74.635 ;
        RECT 108.620 74.600 108.870 74.635 ;
        RECT 109.450 74.600 109.700 74.635 ;
        RECT 110.280 74.600 110.530 74.635 ;
        RECT 111.110 74.600 111.360 74.635 ;
        RECT 111.940 74.625 113.050 74.635 ;
        RECT 64.975 72.575 98.100 74.600 ;
        RECT 98.650 72.575 99.750 74.600 ;
        RECT 100.320 72.575 101.425 74.600 ;
        RECT 101.975 72.575 103.075 74.600 ;
        RECT 103.640 72.575 104.750 74.600 ;
        RECT 105.300 72.575 106.400 74.600 ;
        RECT 106.960 72.575 108.075 74.600 ;
        RECT 108.620 72.575 109.725 74.600 ;
        RECT 110.275 72.575 111.375 74.600 ;
        RECT 64.975 23.400 67.000 72.575 ;
        RECT 97.830 72.530 98.080 72.575 ;
        RECT 98.660 72.530 98.910 72.575 ;
        RECT 99.490 72.530 99.740 72.575 ;
        RECT 100.320 72.530 100.570 72.575 ;
        RECT 101.150 72.530 101.400 72.575 ;
        RECT 101.980 72.530 102.230 72.575 ;
        RECT 102.810 72.530 103.060 72.575 ;
        RECT 103.640 72.530 103.890 72.575 ;
        RECT 104.470 72.530 104.720 72.575 ;
        RECT 105.300 72.530 105.550 72.575 ;
        RECT 106.130 72.530 106.380 72.575 ;
        RECT 106.960 72.530 107.210 72.575 ;
        RECT 107.790 72.530 108.040 72.575 ;
        RECT 108.620 72.530 108.870 72.575 ;
        RECT 109.450 72.530 109.700 72.575 ;
        RECT 110.280 72.530 110.530 72.575 ;
        RECT 111.110 72.530 111.360 72.575 ;
        RECT 111.925 72.550 113.050 74.625 ;
        RECT 113.600 74.600 113.850 74.635 ;
        RECT 114.430 74.600 114.680 74.635 ;
        RECT 115.260 74.600 115.510 74.635 ;
        RECT 116.090 74.600 116.340 74.635 ;
        RECT 116.920 74.600 117.170 74.635 ;
        RECT 117.750 74.600 118.000 74.635 ;
        RECT 118.580 74.600 118.830 74.635 ;
        RECT 119.410 74.600 119.660 74.635 ;
        RECT 120.240 74.600 120.490 74.635 ;
        RECT 121.070 74.600 121.320 74.635 ;
        RECT 121.900 74.600 122.150 74.635 ;
        RECT 122.730 74.600 122.980 74.635 ;
        RECT 123.560 74.600 123.810 74.635 ;
        RECT 124.390 74.600 124.640 74.635 ;
        RECT 125.220 74.600 125.470 74.635 ;
        RECT 126.050 74.600 126.300 74.635 ;
        RECT 126.880 74.600 127.130 74.635 ;
        RECT 127.710 74.600 127.960 74.635 ;
        RECT 128.540 74.600 128.790 74.635 ;
        RECT 129.370 74.600 129.620 74.635 ;
        RECT 130.200 74.600 130.450 74.635 ;
        RECT 131.030 74.600 131.280 74.635 ;
        RECT 131.860 74.600 132.110 74.635 ;
        RECT 132.690 74.600 132.940 74.635 ;
        RECT 133.520 74.600 133.770 74.635 ;
        RECT 134.350 74.600 134.600 74.635 ;
        RECT 135.180 74.600 135.430 74.635 ;
        RECT 136.010 74.600 136.260 74.635 ;
        RECT 136.840 74.600 137.090 74.635 ;
        RECT 137.670 74.600 137.920 74.635 ;
        RECT 138.500 74.600 138.750 74.635 ;
        RECT 139.330 74.600 139.580 74.635 ;
        RECT 140.160 74.600 140.410 74.635 ;
        RECT 140.990 74.600 141.240 74.635 ;
        RECT 141.820 74.600 142.070 74.635 ;
        RECT 142.650 74.600 142.900 74.635 ;
        RECT 143.480 74.600 143.730 74.635 ;
        RECT 144.310 74.600 144.560 74.635 ;
        RECT 145.140 74.600 145.390 74.635 ;
        RECT 145.970 74.600 146.220 74.635 ;
        RECT 146.800 74.600 147.050 74.635 ;
        RECT 147.630 74.600 147.880 74.635 ;
        RECT 148.460 74.600 148.710 74.635 ;
        RECT 149.290 74.600 149.540 74.635 ;
        RECT 150.120 74.600 150.370 74.635 ;
        RECT 150.950 74.600 151.200 74.635 ;
        RECT 151.780 74.600 152.030 74.635 ;
        RECT 152.610 74.600 152.860 74.635 ;
        RECT 153.440 74.600 153.690 74.635 ;
        RECT 154.270 74.600 154.520 74.635 ;
        RECT 155.100 74.600 155.350 74.635 ;
        RECT 155.930 74.600 156.180 74.635 ;
        RECT 156.760 74.600 157.010 74.635 ;
        RECT 157.590 74.600 157.840 74.635 ;
        RECT 158.420 74.600 158.670 74.635 ;
        RECT 159.250 74.600 159.500 74.635 ;
        RECT 160.080 74.600 160.330 74.635 ;
        RECT 160.910 74.600 161.160 74.635 ;
        RECT 161.740 74.600 161.990 74.635 ;
        RECT 162.570 74.600 162.820 74.635 ;
        RECT 163.400 74.600 163.650 74.635 ;
        RECT 164.230 74.600 164.480 74.635 ;
        RECT 165.060 74.600 165.310 74.635 ;
        RECT 165.890 74.600 166.140 74.635 ;
        RECT 166.720 74.600 166.970 74.635 ;
        RECT 167.550 74.600 167.800 74.635 ;
        RECT 168.380 74.600 168.630 74.635 ;
        RECT 169.210 74.600 169.460 74.635 ;
        RECT 170.040 74.600 170.290 74.635 ;
        RECT 170.870 74.600 171.120 74.635 ;
        RECT 171.700 74.600 171.950 74.635 ;
        RECT 172.530 74.600 172.780 74.635 ;
        RECT 173.360 74.600 173.610 74.635 ;
        RECT 174.190 74.600 174.440 74.635 ;
        RECT 175.020 74.600 175.270 74.635 ;
        RECT 175.850 74.600 176.100 74.635 ;
        RECT 176.680 74.600 176.930 74.635 ;
        RECT 177.510 74.600 177.760 74.635 ;
        RECT 178.340 74.600 178.590 74.635 ;
        RECT 179.170 74.600 179.420 74.635 ;
        RECT 113.600 72.575 114.700 74.600 ;
        RECT 115.260 72.575 116.375 74.600 ;
        RECT 116.920 72.575 118.025 74.600 ;
        RECT 118.575 72.575 119.675 74.600 ;
        RECT 120.240 72.575 121.350 74.600 ;
        RECT 121.900 72.575 123.000 74.600 ;
        RECT 123.560 72.575 124.675 74.600 ;
        RECT 125.220 72.575 126.325 74.600 ;
        RECT 126.880 72.575 128.000 74.600 ;
        RECT 128.540 72.575 129.650 74.600 ;
        RECT 130.200 72.575 131.300 74.600 ;
        RECT 131.860 72.575 132.975 74.600 ;
        RECT 133.520 72.575 134.625 74.600 ;
        RECT 135.175 72.575 136.275 74.600 ;
        RECT 136.840 72.575 137.950 74.600 ;
        RECT 138.500 72.575 139.600 74.600 ;
        RECT 140.160 72.575 141.275 74.600 ;
        RECT 141.820 72.575 142.925 74.600 ;
        RECT 143.475 72.575 144.575 74.600 ;
        RECT 145.125 72.575 146.225 74.600 ;
        RECT 146.800 72.575 147.900 74.600 ;
        RECT 148.460 72.575 149.575 74.600 ;
        RECT 150.120 72.575 151.225 74.600 ;
        RECT 151.775 72.575 152.875 74.600 ;
        RECT 153.440 72.575 154.550 74.600 ;
        RECT 155.100 72.575 156.200 74.600 ;
        RECT 156.750 72.575 157.850 74.600 ;
        RECT 158.420 72.575 159.525 74.600 ;
        RECT 160.075 72.575 161.175 74.600 ;
        RECT 161.740 72.575 162.850 74.600 ;
        RECT 163.400 72.575 164.500 74.600 ;
        RECT 165.060 72.575 166.175 74.600 ;
        RECT 166.720 72.575 167.825 74.600 ;
        RECT 168.375 72.575 169.475 74.600 ;
        RECT 170.040 72.575 171.150 74.600 ;
        RECT 171.700 72.575 172.800 74.600 ;
        RECT 173.360 72.575 174.475 74.600 ;
        RECT 175.020 72.575 176.125 74.600 ;
        RECT 176.675 72.575 177.775 74.600 ;
        RECT 178.340 72.575 179.450 74.600 ;
        RECT 111.940 72.530 112.190 72.550 ;
        RECT 112.770 72.530 113.020 72.550 ;
        RECT 113.600 72.530 113.850 72.575 ;
        RECT 114.430 72.530 114.680 72.575 ;
        RECT 115.260 72.530 115.510 72.575 ;
        RECT 116.090 72.530 116.340 72.575 ;
        RECT 116.920 72.530 117.170 72.575 ;
        RECT 117.750 72.530 118.000 72.575 ;
        RECT 118.580 72.530 118.830 72.575 ;
        RECT 119.410 72.530 119.660 72.575 ;
        RECT 120.240 72.530 120.490 72.575 ;
        RECT 121.070 72.530 121.320 72.575 ;
        RECT 121.900 72.530 122.150 72.575 ;
        RECT 122.730 72.530 122.980 72.575 ;
        RECT 123.560 72.530 123.810 72.575 ;
        RECT 124.390 72.530 124.640 72.575 ;
        RECT 125.220 72.530 125.470 72.575 ;
        RECT 126.050 72.530 126.300 72.575 ;
        RECT 126.880 72.530 127.130 72.575 ;
        RECT 127.710 72.530 127.960 72.575 ;
        RECT 128.540 72.530 128.790 72.575 ;
        RECT 129.370 72.530 129.620 72.575 ;
        RECT 130.200 72.530 130.450 72.575 ;
        RECT 131.030 72.530 131.280 72.575 ;
        RECT 131.860 72.530 132.110 72.575 ;
        RECT 132.690 72.530 132.940 72.575 ;
        RECT 133.520 72.530 133.770 72.575 ;
        RECT 134.350 72.530 134.600 72.575 ;
        RECT 135.180 72.530 135.430 72.575 ;
        RECT 136.010 72.530 136.260 72.575 ;
        RECT 136.840 72.530 137.090 72.575 ;
        RECT 137.670 72.530 137.920 72.575 ;
        RECT 138.500 72.530 138.750 72.575 ;
        RECT 139.330 72.530 139.580 72.575 ;
        RECT 140.160 72.530 140.410 72.575 ;
        RECT 140.990 72.530 141.240 72.575 ;
        RECT 141.820 72.530 142.070 72.575 ;
        RECT 142.650 72.530 142.900 72.575 ;
        RECT 143.480 72.530 143.730 72.575 ;
        RECT 144.310 72.530 144.560 72.575 ;
        RECT 145.140 72.530 145.390 72.575 ;
        RECT 145.970 72.530 146.220 72.575 ;
        RECT 146.800 72.530 147.050 72.575 ;
        RECT 147.630 72.530 147.880 72.575 ;
        RECT 148.460 72.530 148.710 72.575 ;
        RECT 149.290 72.530 149.540 72.575 ;
        RECT 150.120 72.530 150.370 72.575 ;
        RECT 150.950 72.530 151.200 72.575 ;
        RECT 151.780 72.530 152.030 72.575 ;
        RECT 152.610 72.530 152.860 72.575 ;
        RECT 153.440 72.530 153.690 72.575 ;
        RECT 154.270 72.530 154.520 72.575 ;
        RECT 155.100 72.530 155.350 72.575 ;
        RECT 155.930 72.530 156.180 72.575 ;
        RECT 156.760 72.530 157.010 72.575 ;
        RECT 157.590 72.530 157.840 72.575 ;
        RECT 158.420 72.530 158.670 72.575 ;
        RECT 159.250 72.530 159.500 72.575 ;
        RECT 160.080 72.530 160.330 72.575 ;
        RECT 160.910 72.530 161.160 72.575 ;
        RECT 161.740 72.530 161.990 72.575 ;
        RECT 162.570 72.530 162.820 72.575 ;
        RECT 163.400 72.530 163.650 72.575 ;
        RECT 164.230 72.530 164.480 72.575 ;
        RECT 165.060 72.530 165.310 72.575 ;
        RECT 165.890 72.530 166.140 72.575 ;
        RECT 166.720 72.530 166.970 72.575 ;
        RECT 167.550 72.530 167.800 72.575 ;
        RECT 168.380 72.530 168.630 72.575 ;
        RECT 169.210 72.530 169.460 72.575 ;
        RECT 170.040 72.530 170.290 72.575 ;
        RECT 170.870 72.530 171.120 72.575 ;
        RECT 171.700 72.530 171.950 72.575 ;
        RECT 172.530 72.530 172.780 72.575 ;
        RECT 173.360 72.530 173.610 72.575 ;
        RECT 174.190 72.530 174.440 72.575 ;
        RECT 175.020 72.530 175.270 72.575 ;
        RECT 175.850 72.530 176.100 72.575 ;
        RECT 176.680 72.530 176.930 72.575 ;
        RECT 177.510 72.530 177.760 72.575 ;
        RECT 178.340 72.530 178.590 72.575 ;
        RECT 179.170 72.530 179.420 72.575 ;
        RECT 179.900 72.525 180.350 74.650 ;
        RECT 180.650 72.525 181.250 74.650 ;
        RECT 181.660 74.600 181.910 74.635 ;
        RECT 182.490 74.600 182.740 74.635 ;
        RECT 183.320 74.600 183.570 74.635 ;
        RECT 184.150 74.600 184.400 74.635 ;
        RECT 184.980 74.600 185.230 74.635 ;
        RECT 185.810 74.600 186.060 74.635 ;
        RECT 186.640 74.600 186.890 74.635 ;
        RECT 187.470 74.600 187.720 74.635 ;
        RECT 188.300 74.600 188.550 74.635 ;
        RECT 189.130 74.600 189.380 74.635 ;
        RECT 189.960 74.600 190.210 74.635 ;
        RECT 190.790 74.600 191.040 74.635 ;
        RECT 191.620 74.600 191.870 74.635 ;
        RECT 192.450 74.600 192.700 74.635 ;
        RECT 193.280 74.600 193.530 74.635 ;
        RECT 194.110 74.600 194.360 74.635 ;
        RECT 194.940 74.600 195.190 74.635 ;
        RECT 195.770 74.600 196.020 74.635 ;
        RECT 196.600 74.600 196.850 74.635 ;
        RECT 197.430 74.600 197.680 74.635 ;
        RECT 198.260 74.600 198.510 74.635 ;
        RECT 199.090 74.600 199.340 74.635 ;
        RECT 199.920 74.600 200.170 74.635 ;
        RECT 200.750 74.600 201.000 74.635 ;
        RECT 201.580 74.600 201.830 74.635 ;
        RECT 202.410 74.600 202.660 74.635 ;
        RECT 203.240 74.600 203.490 74.635 ;
        RECT 204.070 74.600 204.320 74.635 ;
        RECT 204.900 74.600 205.150 74.635 ;
        RECT 205.730 74.600 205.980 74.635 ;
        RECT 206.560 74.600 206.810 74.635 ;
        RECT 207.390 74.600 207.640 74.635 ;
        RECT 208.220 74.600 208.470 74.635 ;
        RECT 209.050 74.600 209.300 74.635 ;
        RECT 209.880 74.600 210.130 74.635 ;
        RECT 210.710 74.600 210.960 74.635 ;
        RECT 211.540 74.600 211.790 74.635 ;
        RECT 181.660 72.575 182.775 74.600 ;
        RECT 183.320 72.575 184.425 74.600 ;
        RECT 184.975 72.575 186.075 74.600 ;
        RECT 186.640 72.575 187.750 74.600 ;
        RECT 188.300 72.575 189.400 74.600 ;
        RECT 189.960 72.575 191.075 74.600 ;
        RECT 191.620 72.575 192.725 74.600 ;
        RECT 193.275 72.575 194.375 74.600 ;
        RECT 194.940 72.575 196.050 74.600 ;
        RECT 196.600 72.575 197.700 74.600 ;
        RECT 198.260 72.575 199.375 74.600 ;
        RECT 199.920 72.575 201.025 74.600 ;
        RECT 201.575 72.575 202.675 74.600 ;
        RECT 203.240 72.575 204.350 74.600 ;
        RECT 204.900 72.575 206.000 74.600 ;
        RECT 206.560 72.575 207.675 74.600 ;
        RECT 208.220 72.575 209.325 74.600 ;
        RECT 209.875 72.575 210.975 74.600 ;
        RECT 211.540 72.575 214.125 74.600 ;
        RECT 181.660 72.530 181.910 72.575 ;
        RECT 182.490 72.530 182.740 72.575 ;
        RECT 183.320 72.530 183.570 72.575 ;
        RECT 184.150 72.530 184.400 72.575 ;
        RECT 184.980 72.530 185.230 72.575 ;
        RECT 185.810 72.530 186.060 72.575 ;
        RECT 186.640 72.530 186.890 72.575 ;
        RECT 187.470 72.530 187.720 72.575 ;
        RECT 188.300 72.530 188.550 72.575 ;
        RECT 189.130 72.530 189.380 72.575 ;
        RECT 189.960 72.530 190.210 72.575 ;
        RECT 190.790 72.530 191.040 72.575 ;
        RECT 191.620 72.530 191.870 72.575 ;
        RECT 192.450 72.530 192.700 72.575 ;
        RECT 193.280 72.530 193.530 72.575 ;
        RECT 194.110 72.530 194.360 72.575 ;
        RECT 194.940 72.530 195.190 72.575 ;
        RECT 195.770 72.530 196.020 72.575 ;
        RECT 196.600 72.530 196.850 72.575 ;
        RECT 197.430 72.530 197.680 72.575 ;
        RECT 198.260 72.530 198.510 72.575 ;
        RECT 199.090 72.530 199.340 72.575 ;
        RECT 199.920 72.530 200.170 72.575 ;
        RECT 200.750 72.530 201.000 72.575 ;
        RECT 201.580 72.530 201.830 72.575 ;
        RECT 202.410 72.530 202.660 72.575 ;
        RECT 203.240 72.530 203.490 72.575 ;
        RECT 204.070 72.530 204.320 72.575 ;
        RECT 204.900 72.530 205.150 72.575 ;
        RECT 205.730 72.530 205.980 72.575 ;
        RECT 206.560 72.530 206.810 72.575 ;
        RECT 207.390 72.530 207.640 72.575 ;
        RECT 208.220 72.530 208.470 72.575 ;
        RECT 209.050 72.530 209.300 72.575 ;
        RECT 209.880 72.530 210.130 72.575 ;
        RECT 210.710 72.530 210.960 72.575 ;
        RECT 211.540 72.530 211.790 72.575 ;
        RECT 215.625 71.900 228.050 75.945 ;
        RECT 75.275 68.025 97.300 71.900 ;
        RECT 97.830 70.600 98.080 70.640 ;
        RECT 98.660 70.600 98.910 70.640 ;
        RECT 99.490 70.600 99.740 70.640 ;
        RECT 100.320 70.600 100.570 70.640 ;
        RECT 101.150 70.600 101.400 70.640 ;
        RECT 101.980 70.600 102.230 70.640 ;
        RECT 102.810 70.600 103.060 70.640 ;
        RECT 103.640 70.600 103.890 70.640 ;
        RECT 104.470 70.600 104.720 70.640 ;
        RECT 105.300 70.600 105.550 70.640 ;
        RECT 106.130 70.600 106.380 70.640 ;
        RECT 106.960 70.600 107.210 70.640 ;
        RECT 107.790 70.600 108.040 70.640 ;
        RECT 108.620 70.600 108.870 70.640 ;
        RECT 109.450 70.600 109.700 70.640 ;
        RECT 110.280 70.600 110.530 70.640 ;
        RECT 111.110 70.600 111.360 70.640 ;
        RECT 111.940 70.600 112.190 70.640 ;
        RECT 112.770 70.600 113.020 70.640 ;
        RECT 113.600 70.600 113.850 70.640 ;
        RECT 114.430 70.600 114.680 70.640 ;
        RECT 115.260 70.600 115.510 70.640 ;
        RECT 116.090 70.600 116.340 70.640 ;
        RECT 116.920 70.600 117.170 70.640 ;
        RECT 117.750 70.600 118.000 70.640 ;
        RECT 118.580 70.600 118.830 70.640 ;
        RECT 119.410 70.600 119.660 70.640 ;
        RECT 120.240 70.600 120.490 70.640 ;
        RECT 121.070 70.600 121.320 70.640 ;
        RECT 121.900 70.600 122.150 70.640 ;
        RECT 122.730 70.600 122.980 70.640 ;
        RECT 123.560 70.600 123.810 70.640 ;
        RECT 124.390 70.600 124.640 70.640 ;
        RECT 125.220 70.600 125.470 70.640 ;
        RECT 126.050 70.600 126.300 70.640 ;
        RECT 126.880 70.600 127.130 70.640 ;
        RECT 97.825 68.575 98.925 70.600 ;
        RECT 99.475 68.575 100.600 70.600 ;
        RECT 101.150 68.575 102.250 70.600 ;
        RECT 102.800 68.575 103.900 70.600 ;
        RECT 104.470 68.575 105.575 70.600 ;
        RECT 106.125 68.575 107.225 70.600 ;
        RECT 107.775 68.575 108.875 70.600 ;
        RECT 109.450 68.575 110.550 70.600 ;
        RECT 111.100 68.575 112.200 70.600 ;
        RECT 112.770 68.575 113.875 70.600 ;
        RECT 114.425 68.575 115.525 70.600 ;
        RECT 116.090 68.575 117.200 70.600 ;
        RECT 117.750 68.575 118.850 70.600 ;
        RECT 119.400 68.575 120.500 70.600 ;
        RECT 121.070 68.575 122.175 70.600 ;
        RECT 122.725 68.575 123.825 70.600 ;
        RECT 124.390 68.575 125.500 70.600 ;
        RECT 126.050 68.575 127.150 70.600 ;
        RECT 97.830 68.535 98.080 68.575 ;
        RECT 98.660 68.535 98.910 68.575 ;
        RECT 99.490 68.535 99.740 68.575 ;
        RECT 100.320 68.535 100.570 68.575 ;
        RECT 101.150 68.535 101.400 68.575 ;
        RECT 101.980 68.535 102.230 68.575 ;
        RECT 102.810 68.535 103.060 68.575 ;
        RECT 103.640 68.535 103.890 68.575 ;
        RECT 104.470 68.535 104.720 68.575 ;
        RECT 105.300 68.535 105.550 68.575 ;
        RECT 106.130 68.535 106.380 68.575 ;
        RECT 106.960 68.535 107.210 68.575 ;
        RECT 107.790 68.535 108.040 68.575 ;
        RECT 108.620 68.535 108.870 68.575 ;
        RECT 109.450 68.535 109.700 68.575 ;
        RECT 110.280 68.535 110.530 68.575 ;
        RECT 111.110 68.535 111.360 68.575 ;
        RECT 111.940 68.535 112.190 68.575 ;
        RECT 112.770 68.535 113.020 68.575 ;
        RECT 113.600 68.535 113.850 68.575 ;
        RECT 114.430 68.535 114.680 68.575 ;
        RECT 115.260 68.535 115.510 68.575 ;
        RECT 116.090 68.535 116.340 68.575 ;
        RECT 116.920 68.535 117.170 68.575 ;
        RECT 117.750 68.535 118.000 68.575 ;
        RECT 118.580 68.535 118.830 68.575 ;
        RECT 119.410 68.535 119.660 68.575 ;
        RECT 120.240 68.535 120.490 68.575 ;
        RECT 121.070 68.535 121.320 68.575 ;
        RECT 121.900 68.535 122.150 68.575 ;
        RECT 122.730 68.535 122.980 68.575 ;
        RECT 123.560 68.535 123.810 68.575 ;
        RECT 124.390 68.535 124.640 68.575 ;
        RECT 125.220 68.535 125.470 68.575 ;
        RECT 126.050 68.535 126.300 68.575 ;
        RECT 126.880 68.535 127.130 68.575 ;
        RECT 127.675 68.525 128.825 70.650 ;
        RECT 129.370 70.600 129.620 70.640 ;
        RECT 130.200 70.600 130.450 70.640 ;
        RECT 131.030 70.600 131.280 70.640 ;
        RECT 131.860 70.600 132.110 70.640 ;
        RECT 132.690 70.600 132.940 70.640 ;
        RECT 133.520 70.600 133.770 70.640 ;
        RECT 134.350 70.600 134.600 70.640 ;
        RECT 135.180 70.600 135.430 70.640 ;
        RECT 136.010 70.600 136.260 70.640 ;
        RECT 136.840 70.600 137.090 70.640 ;
        RECT 137.670 70.600 137.920 70.640 ;
        RECT 138.500 70.600 138.750 70.640 ;
        RECT 139.330 70.600 139.580 70.640 ;
        RECT 140.160 70.600 140.410 70.640 ;
        RECT 140.990 70.600 141.240 70.640 ;
        RECT 141.820 70.600 142.070 70.640 ;
        RECT 142.650 70.600 142.900 70.640 ;
        RECT 143.480 70.600 143.730 70.640 ;
        RECT 144.310 70.600 144.560 70.640 ;
        RECT 145.140 70.600 145.390 70.640 ;
        RECT 145.970 70.600 146.220 70.640 ;
        RECT 146.800 70.600 147.050 70.640 ;
        RECT 147.630 70.600 147.880 70.640 ;
        RECT 148.460 70.600 148.710 70.640 ;
        RECT 149.290 70.600 149.540 70.640 ;
        RECT 150.120 70.600 150.370 70.640 ;
        RECT 150.950 70.600 151.200 70.640 ;
        RECT 151.780 70.600 152.030 70.640 ;
        RECT 152.610 70.600 152.860 70.640 ;
        RECT 153.440 70.600 153.690 70.640 ;
        RECT 154.270 70.600 154.520 70.640 ;
        RECT 155.100 70.600 155.350 70.640 ;
        RECT 155.930 70.600 156.180 70.640 ;
        RECT 156.760 70.600 157.010 70.640 ;
        RECT 157.590 70.600 157.840 70.640 ;
        RECT 158.420 70.600 158.670 70.640 ;
        RECT 159.250 70.600 159.500 70.640 ;
        RECT 160.080 70.600 160.330 70.640 ;
        RECT 160.910 70.600 161.160 70.640 ;
        RECT 161.740 70.600 161.990 70.640 ;
        RECT 162.570 70.600 162.820 70.640 ;
        RECT 163.400 70.600 163.650 70.640 ;
        RECT 164.230 70.600 164.480 70.640 ;
        RECT 165.060 70.600 165.310 70.640 ;
        RECT 165.890 70.600 166.140 70.640 ;
        RECT 166.720 70.600 166.970 70.640 ;
        RECT 167.550 70.600 167.800 70.640 ;
        RECT 168.380 70.600 168.630 70.640 ;
        RECT 169.210 70.600 169.460 70.640 ;
        RECT 170.040 70.600 170.290 70.640 ;
        RECT 170.870 70.600 171.120 70.640 ;
        RECT 171.700 70.600 171.950 70.640 ;
        RECT 172.530 70.600 172.780 70.640 ;
        RECT 173.360 70.600 173.610 70.640 ;
        RECT 174.190 70.600 174.440 70.640 ;
        RECT 175.020 70.600 175.270 70.640 ;
        RECT 175.850 70.600 176.100 70.640 ;
        RECT 176.680 70.600 176.930 70.640 ;
        RECT 177.510 70.600 177.760 70.640 ;
        RECT 178.340 70.600 178.590 70.640 ;
        RECT 179.170 70.600 179.420 70.640 ;
        RECT 180.000 70.600 180.250 70.640 ;
        RECT 180.830 70.600 181.080 70.640 ;
        RECT 181.660 70.600 181.910 70.640 ;
        RECT 182.490 70.600 182.740 70.640 ;
        RECT 183.320 70.600 183.570 70.640 ;
        RECT 184.150 70.600 184.400 70.640 ;
        RECT 184.980 70.600 185.230 70.640 ;
        RECT 185.810 70.600 186.060 70.640 ;
        RECT 186.640 70.600 186.890 70.640 ;
        RECT 187.470 70.600 187.720 70.640 ;
        RECT 188.300 70.600 188.550 70.640 ;
        RECT 189.130 70.600 189.380 70.640 ;
        RECT 189.960 70.600 190.210 70.640 ;
        RECT 190.790 70.600 191.040 70.640 ;
        RECT 191.620 70.600 191.870 70.640 ;
        RECT 192.450 70.600 192.700 70.640 ;
        RECT 193.280 70.600 193.530 70.640 ;
        RECT 194.110 70.600 194.360 70.640 ;
        RECT 194.940 70.600 195.190 70.640 ;
        RECT 195.770 70.600 196.020 70.640 ;
        RECT 196.600 70.600 196.850 70.640 ;
        RECT 197.430 70.600 197.680 70.640 ;
        RECT 198.260 70.600 198.510 70.640 ;
        RECT 199.090 70.600 199.340 70.640 ;
        RECT 199.920 70.600 200.170 70.640 ;
        RECT 200.750 70.600 201.000 70.640 ;
        RECT 201.580 70.600 201.830 70.640 ;
        RECT 202.410 70.600 202.660 70.640 ;
        RECT 203.240 70.600 203.490 70.640 ;
        RECT 204.070 70.600 204.320 70.640 ;
        RECT 204.900 70.600 205.150 70.640 ;
        RECT 205.730 70.600 205.980 70.640 ;
        RECT 206.560 70.600 206.810 70.640 ;
        RECT 207.390 70.600 207.640 70.640 ;
        RECT 208.220 70.600 208.470 70.640 ;
        RECT 209.050 70.600 209.300 70.640 ;
        RECT 209.880 70.600 210.130 70.640 ;
        RECT 210.710 70.600 210.960 70.640 ;
        RECT 211.540 70.600 211.790 70.640 ;
        RECT 129.370 68.575 130.475 70.600 ;
        RECT 131.025 68.575 132.125 70.600 ;
        RECT 132.690 68.575 133.800 70.600 ;
        RECT 134.350 68.575 135.450 70.600 ;
        RECT 136.000 68.575 137.100 70.600 ;
        RECT 137.670 68.575 138.775 70.600 ;
        RECT 139.325 68.575 140.425 70.600 ;
        RECT 140.990 68.575 142.100 70.600 ;
        RECT 142.650 68.575 143.750 70.600 ;
        RECT 144.310 68.575 145.425 70.600 ;
        RECT 145.970 68.575 147.075 70.600 ;
        RECT 147.625 68.575 148.725 70.600 ;
        RECT 149.290 68.575 150.400 70.600 ;
        RECT 150.950 68.575 152.050 70.600 ;
        RECT 152.610 68.575 153.725 70.600 ;
        RECT 154.270 68.575 155.375 70.600 ;
        RECT 155.925 68.575 157.025 70.600 ;
        RECT 157.590 68.575 158.700 70.600 ;
        RECT 159.250 68.575 160.350 70.600 ;
        RECT 160.900 68.575 162.000 70.600 ;
        RECT 162.570 68.575 163.675 70.600 ;
        RECT 164.225 68.575 165.325 70.600 ;
        RECT 165.890 68.575 167.000 70.600 ;
        RECT 167.550 68.575 168.650 70.600 ;
        RECT 169.200 68.575 170.300 70.600 ;
        RECT 170.850 68.575 171.950 70.600 ;
        RECT 172.525 68.575 173.625 70.600 ;
        RECT 174.190 68.575 175.300 70.600 ;
        RECT 175.850 68.575 176.950 70.600 ;
        RECT 177.500 68.575 178.600 70.600 ;
        RECT 179.170 68.575 180.275 70.600 ;
        RECT 180.825 68.575 181.925 70.600 ;
        RECT 182.490 68.575 183.600 70.600 ;
        RECT 184.150 68.575 185.250 70.600 ;
        RECT 185.810 68.575 186.925 70.600 ;
        RECT 187.470 68.575 188.575 70.600 ;
        RECT 189.125 68.575 190.225 70.600 ;
        RECT 190.775 68.575 191.875 70.600 ;
        RECT 192.450 68.575 193.550 70.600 ;
        RECT 194.100 68.575 195.200 70.600 ;
        RECT 195.750 68.575 196.850 70.600 ;
        RECT 197.425 68.575 198.525 70.600 ;
        RECT 199.090 68.575 200.200 70.600 ;
        RECT 200.750 68.575 201.850 70.600 ;
        RECT 202.400 68.575 203.500 70.600 ;
        RECT 204.070 68.575 205.175 70.600 ;
        RECT 205.725 68.575 206.825 70.600 ;
        RECT 207.375 68.575 208.475 70.600 ;
        RECT 209.050 68.575 210.150 70.600 ;
        RECT 210.700 68.575 211.800 70.600 ;
        RECT 212.325 68.850 228.050 71.900 ;
        RECT 230.000 79.625 230.600 86.300 ;
        RECT 231.050 84.645 266.400 85.500 ;
        RECT 231.045 84.300 266.400 84.645 ;
        RECT 231.045 84.295 234.650 84.300 ;
        RECT 235.645 84.295 248.450 84.300 ;
        RECT 231.050 84.275 234.650 84.295 ;
        RECT 231.050 83.550 232.050 84.275 ;
        RECT 233.650 84.095 234.650 84.275 ;
        RECT 233.645 83.770 234.650 84.095 ;
        RECT 233.650 83.550 234.650 83.770 ;
        RECT 231.050 83.545 232.275 83.550 ;
        RECT 231.050 80.550 232.480 83.545 ;
        RECT 232.675 80.550 233.025 83.550 ;
        RECT 233.425 83.545 234.650 83.550 ;
        RECT 233.210 80.550 234.650 83.545 ;
        RECT 235.650 84.275 248.450 84.295 ;
        RECT 235.650 83.550 236.650 84.275 ;
        RECT 238.250 84.095 241.525 84.275 ;
        RECT 242.575 84.095 245.850 84.275 ;
        RECT 247.450 84.095 248.450 84.275 ;
        RECT 238.245 83.775 241.525 84.095 ;
        RECT 238.245 83.770 241.250 83.775 ;
        RECT 242.570 83.770 245.850 84.095 ;
        RECT 247.445 83.770 248.450 84.095 ;
        RECT 238.250 83.550 241.250 83.770 ;
        RECT 242.850 83.550 245.850 83.770 ;
        RECT 247.450 83.550 248.450 83.770 ;
        RECT 235.650 83.545 236.875 83.550 ;
        RECT 235.650 80.550 237.080 83.545 ;
        RECT 237.275 80.550 237.625 83.550 ;
        RECT 238.025 83.545 241.475 83.550 ;
        RECT 237.810 80.550 241.680 83.545 ;
        RECT 241.875 80.550 242.225 83.550 ;
        RECT 242.625 83.545 246.075 83.550 ;
        RECT 242.410 80.550 246.280 83.545 ;
        RECT 246.475 80.550 246.825 83.550 ;
        RECT 247.225 83.545 248.450 83.550 ;
        RECT 247.010 80.550 248.450 83.545 ;
        RECT 249.450 84.100 250.450 84.300 ;
        RECT 249.450 83.775 250.455 84.100 ;
        RECT 249.450 83.550 250.450 83.775 ;
        RECT 249.450 80.550 250.880 83.550 ;
        RECT 251.075 80.550 251.400 83.550 ;
        RECT 251.600 80.550 251.850 84.300 ;
        RECT 252.050 80.550 252.375 83.550 ;
        RECT 252.550 80.550 252.800 84.300 ;
        RECT 253.950 84.150 266.400 84.300 ;
        RECT 253.950 83.550 254.950 84.150 ;
        RECT 253.000 80.550 253.325 83.550 ;
        RECT 253.530 80.550 254.950 83.550 ;
        RECT 231.770 80.545 232.000 80.550 ;
        RECT 232.250 80.545 232.480 80.550 ;
        RECT 232.730 80.545 232.960 80.550 ;
        RECT 233.210 80.545 233.440 80.550 ;
        RECT 233.690 80.545 233.920 80.550 ;
        RECT 236.370 80.545 236.600 80.550 ;
        RECT 236.850 80.545 237.080 80.550 ;
        RECT 237.330 80.545 237.560 80.550 ;
        RECT 237.810 80.545 238.040 80.550 ;
        RECT 238.290 80.545 238.520 80.550 ;
        RECT 240.970 80.545 241.200 80.550 ;
        RECT 241.450 80.545 241.680 80.550 ;
        RECT 241.930 80.545 242.160 80.550 ;
        RECT 242.410 80.545 242.640 80.550 ;
        RECT 242.890 80.545 243.120 80.550 ;
        RECT 245.570 80.545 245.800 80.550 ;
        RECT 246.050 80.545 246.280 80.550 ;
        RECT 246.530 80.545 246.760 80.550 ;
        RECT 247.010 80.545 247.240 80.550 ;
        RECT 247.490 80.545 247.720 80.550 ;
        RECT 232.450 80.345 233.250 80.350 ;
        RECT 237.050 80.345 237.850 80.350 ;
        RECT 242.100 80.345 242.475 80.350 ;
        RECT 246.250 80.345 247.050 80.350 ;
        RECT 232.445 79.970 233.250 80.345 ;
        RECT 237.045 79.970 237.850 80.345 ;
        RECT 242.095 79.970 242.475 80.345 ;
        RECT 246.245 79.970 247.050 80.345 ;
        RECT 232.450 79.625 233.250 79.970 ;
        RECT 237.050 79.625 237.850 79.970 ;
        RECT 242.100 79.625 242.475 79.970 ;
        RECT 246.250 79.625 247.050 79.970 ;
        RECT 250.825 79.975 253.580 80.350 ;
        RECT 250.825 79.625 253.575 79.975 ;
        RECT 230.000 79.025 233.250 79.625 ;
        RECT 234.900 79.025 237.850 79.625 ;
        RECT 239.500 79.025 242.475 79.625 ;
        RECT 244.775 79.025 247.050 79.625 ;
        RECT 248.700 79.025 253.575 79.625 ;
        RECT 230.000 70.325 230.600 79.025 ;
        RECT 232.450 78.350 233.250 79.025 ;
        RECT 237.050 78.350 237.850 79.025 ;
        RECT 242.100 78.350 242.475 79.025 ;
        RECT 246.250 78.350 247.050 79.025 ;
        RECT 250.825 78.675 253.575 79.025 ;
        RECT 250.825 78.350 253.580 78.675 ;
        RECT 256.625 78.600 271.250 78.950 ;
        RECT 231.050 77.150 232.485 78.150 ;
        RECT 232.675 77.150 233.025 78.150 ;
        RECT 233.215 77.150 237.085 78.150 ;
        RECT 237.275 77.150 237.625 78.150 ;
        RECT 237.815 77.150 239.250 78.150 ;
        RECT 231.050 76.450 232.050 77.150 ;
        RECT 233.650 76.450 236.650 77.150 ;
        RECT 238.250 76.450 239.250 77.150 ;
        RECT 240.250 77.150 241.685 78.150 ;
        RECT 241.875 77.150 242.225 78.150 ;
        RECT 242.415 77.150 243.850 78.150 ;
        RECT 240.250 76.950 241.250 77.150 ;
        RECT 242.850 76.950 243.850 77.150 ;
        RECT 240.250 76.450 241.525 76.950 ;
        RECT 242.575 76.450 243.850 76.950 ;
        RECT 244.850 77.150 246.285 78.150 ;
        RECT 246.475 77.150 246.825 78.150 ;
        RECT 247.015 77.150 250.880 78.150 ;
        RECT 251.075 77.150 251.400 78.150 ;
        RECT 244.850 76.450 245.850 77.150 ;
        RECT 247.450 77.125 250.880 77.150 ;
        RECT 247.450 76.450 250.875 77.125 ;
        RECT 251.600 76.450 251.850 78.150 ;
        RECT 252.050 77.150 252.375 78.150 ;
        RECT 252.550 76.450 252.800 78.150 ;
        RECT 253.000 77.150 253.325 78.150 ;
        RECT 253.525 76.450 254.950 78.150 ;
        RECT 256.625 78.050 271.250 78.425 ;
        RECT 231.050 76.100 254.955 76.450 ;
        RECT 231.050 75.350 233.700 75.355 ;
        RECT 231.050 75.000 254.955 75.350 ;
        RECT 231.050 71.250 231.425 75.000 ;
        RECT 231.950 74.450 232.800 74.830 ;
        RECT 231.775 70.325 232.025 74.275 ;
        RECT 232.200 71.250 232.550 74.275 ;
        RECT 232.725 70.325 232.975 74.275 ;
        RECT 233.325 71.250 233.700 75.000 ;
        RECT 235.645 74.995 248.450 75.000 ;
        RECT 235.650 74.975 248.450 74.995 ;
        RECT 235.650 74.250 236.650 74.975 ;
        RECT 238.250 74.795 241.525 74.975 ;
        RECT 242.575 74.795 245.850 74.975 ;
        RECT 247.450 74.795 248.450 74.975 ;
        RECT 238.245 74.475 241.525 74.795 ;
        RECT 238.245 74.470 241.250 74.475 ;
        RECT 242.570 74.470 245.850 74.795 ;
        RECT 247.445 74.470 248.450 74.795 ;
        RECT 238.250 74.250 241.250 74.470 ;
        RECT 242.850 74.250 245.850 74.470 ;
        RECT 247.450 74.250 248.450 74.470 ;
        RECT 235.650 74.245 236.875 74.250 ;
        RECT 235.650 71.250 237.080 74.245 ;
        RECT 237.275 71.250 237.625 74.250 ;
        RECT 238.025 74.245 241.475 74.250 ;
        RECT 237.810 71.250 241.680 74.245 ;
        RECT 241.875 71.250 242.225 74.250 ;
        RECT 242.625 74.245 246.075 74.250 ;
        RECT 242.410 71.250 246.280 74.245 ;
        RECT 246.475 71.250 246.825 74.250 ;
        RECT 247.225 74.245 248.450 74.250 ;
        RECT 247.010 71.250 248.450 74.245 ;
        RECT 249.450 74.800 250.450 75.000 ;
        RECT 249.450 74.475 250.455 74.800 ;
        RECT 249.450 74.250 250.450 74.475 ;
        RECT 249.450 71.250 250.880 74.250 ;
        RECT 251.075 71.250 251.400 74.250 ;
        RECT 251.600 71.250 251.850 75.000 ;
        RECT 252.050 71.250 252.375 74.250 ;
        RECT 252.550 71.250 252.800 75.000 ;
        RECT 253.950 74.250 254.950 75.000 ;
        RECT 253.000 71.250 253.325 74.250 ;
        RECT 253.530 71.250 254.950 74.250 ;
        RECT 256.625 71.250 256.975 78.050 ;
        RECT 257.540 78.045 259.290 78.050 ;
        RECT 268.590 78.045 270.340 78.050 ;
        RECT 257.345 77.775 257.575 77.845 ;
        RECT 257.825 77.775 258.055 77.845 ;
        RECT 258.305 77.775 258.535 77.845 ;
        RECT 258.785 77.775 259.015 77.845 ;
        RECT 259.265 77.775 259.495 77.845 ;
        RECT 259.745 77.775 259.975 77.845 ;
        RECT 257.300 76.600 259.500 77.775 ;
        RECT 259.700 76.600 260.025 77.775 ;
        RECT 257.345 74.845 257.575 76.600 ;
        RECT 257.825 74.845 258.055 76.600 ;
        RECT 258.305 74.845 258.535 76.600 ;
        RECT 258.785 74.845 259.015 76.600 ;
        RECT 259.225 76.575 259.500 76.600 ;
        RECT 259.225 74.850 259.550 76.575 ;
        RECT 259.265 74.845 259.495 74.850 ;
        RECT 259.745 74.845 259.975 76.600 ;
        RECT 260.225 76.025 260.455 77.845 ;
        RECT 260.705 77.775 260.935 77.845 ;
        RECT 260.650 76.600 260.975 77.775 ;
        RECT 260.175 74.850 260.500 76.025 ;
        RECT 260.225 74.845 260.455 74.850 ;
        RECT 260.705 74.845 260.935 76.600 ;
        RECT 261.185 76.025 261.415 77.845 ;
        RECT 261.665 77.775 261.895 77.845 ;
        RECT 261.625 76.600 261.950 77.775 ;
        RECT 261.125 74.850 261.475 76.025 ;
        RECT 261.185 74.845 261.415 74.850 ;
        RECT 261.665 74.845 261.895 76.600 ;
        RECT 262.145 76.025 262.375 77.845 ;
        RECT 262.625 77.775 262.855 77.845 ;
        RECT 262.575 76.600 262.900 77.775 ;
        RECT 262.100 74.850 262.425 76.025 ;
        RECT 262.145 74.845 262.375 74.850 ;
        RECT 262.625 74.845 262.855 76.600 ;
        RECT 263.105 76.025 263.335 77.845 ;
        RECT 263.585 77.775 263.815 77.845 ;
        RECT 263.525 76.600 263.875 77.775 ;
        RECT 263.050 74.850 263.375 76.025 ;
        RECT 263.105 74.845 263.335 74.850 ;
        RECT 263.585 74.845 263.815 76.600 ;
        RECT 264.065 76.025 264.295 77.845 ;
        RECT 264.545 77.775 264.775 77.845 ;
        RECT 264.500 76.600 264.825 77.775 ;
        RECT 264.025 74.850 264.350 76.025 ;
        RECT 264.065 74.845 264.295 74.850 ;
        RECT 264.545 74.845 264.775 76.600 ;
        RECT 265.025 76.025 265.255 77.845 ;
        RECT 265.505 77.775 265.735 77.845 ;
        RECT 265.450 76.600 265.775 77.775 ;
        RECT 264.975 74.850 265.300 76.025 ;
        RECT 265.025 74.845 265.255 74.850 ;
        RECT 265.505 74.845 265.735 76.600 ;
        RECT 265.985 76.025 266.215 77.845 ;
        RECT 266.465 77.775 266.695 77.845 ;
        RECT 266.425 76.600 266.750 77.775 ;
        RECT 265.925 74.850 266.250 76.025 ;
        RECT 265.985 74.845 266.215 74.850 ;
        RECT 266.465 74.845 266.695 76.600 ;
        RECT 266.945 76.025 267.175 77.845 ;
        RECT 267.425 77.775 267.655 77.845 ;
        RECT 267.375 76.600 267.700 77.775 ;
        RECT 266.900 74.850 267.225 76.025 ;
        RECT 266.945 74.845 267.175 74.850 ;
        RECT 267.425 74.845 267.655 76.600 ;
        RECT 267.905 76.025 268.135 77.845 ;
        RECT 268.385 77.775 268.615 77.845 ;
        RECT 268.865 77.775 269.095 77.845 ;
        RECT 269.345 77.775 269.575 77.845 ;
        RECT 269.825 77.775 270.055 77.845 ;
        RECT 270.305 77.775 270.535 77.845 ;
        RECT 268.325 76.600 270.575 77.775 ;
        RECT 267.850 74.850 268.175 76.025 ;
        RECT 267.905 74.845 268.135 74.850 ;
        RECT 268.385 74.845 268.615 76.600 ;
        RECT 268.865 74.845 269.095 76.600 ;
        RECT 269.345 74.845 269.575 76.600 ;
        RECT 269.825 74.845 270.055 76.600 ;
        RECT 270.305 74.845 270.535 76.600 ;
        RECT 257.525 72.650 270.350 74.650 ;
        RECT 257.345 71.800 257.575 72.450 ;
        RECT 257.825 71.800 258.055 72.450 ;
        RECT 258.305 71.800 258.535 72.450 ;
        RECT 258.785 71.800 259.015 72.450 ;
        RECT 259.225 71.825 259.550 72.450 ;
        RECT 259.225 71.800 259.525 71.825 ;
        RECT 259.745 71.800 259.975 72.450 ;
        RECT 260.175 72.050 260.500 72.450 ;
        RECT 257.300 71.400 259.525 71.800 ;
        RECT 259.700 71.400 260.025 71.800 ;
        RECT 260.225 71.450 260.455 72.050 ;
        RECT 260.705 71.800 260.935 72.450 ;
        RECT 261.125 72.050 261.475 72.450 ;
        RECT 260.650 71.400 261.000 71.800 ;
        RECT 261.185 71.450 261.415 72.050 ;
        RECT 261.665 71.800 261.895 72.450 ;
        RECT 262.100 72.050 262.425 72.450 ;
        RECT 261.625 71.400 261.950 71.800 ;
        RECT 262.145 71.450 262.375 72.050 ;
        RECT 262.625 71.800 262.855 72.450 ;
        RECT 263.050 72.050 263.375 72.450 ;
        RECT 262.575 71.400 262.900 71.800 ;
        RECT 263.105 71.450 263.335 72.050 ;
        RECT 263.585 71.800 263.815 72.450 ;
        RECT 264.025 72.050 264.350 72.450 ;
        RECT 263.525 71.400 263.875 71.800 ;
        RECT 264.065 71.450 264.295 72.050 ;
        RECT 264.545 71.800 264.775 72.450 ;
        RECT 264.975 72.050 265.300 72.450 ;
        RECT 264.500 71.400 264.825 71.800 ;
        RECT 265.025 71.450 265.255 72.050 ;
        RECT 265.505 71.800 265.735 72.450 ;
        RECT 265.925 72.050 266.275 72.450 ;
        RECT 265.450 71.400 265.800 71.800 ;
        RECT 265.985 71.450 266.215 72.050 ;
        RECT 266.465 71.800 266.695 72.450 ;
        RECT 266.900 72.050 267.225 72.450 ;
        RECT 266.425 71.400 266.750 71.800 ;
        RECT 266.945 71.450 267.175 72.050 ;
        RECT 267.425 71.800 267.655 72.450 ;
        RECT 267.850 72.050 268.200 72.450 ;
        RECT 267.375 71.400 267.700 71.800 ;
        RECT 267.905 71.450 268.135 72.050 ;
        RECT 268.385 71.800 268.615 72.450 ;
        RECT 268.865 71.800 269.095 72.450 ;
        RECT 269.345 71.800 269.575 72.450 ;
        RECT 269.825 71.800 270.055 72.450 ;
        RECT 270.305 71.800 270.535 72.450 ;
        RECT 268.325 71.400 270.575 71.800 ;
        RECT 270.900 71.250 271.250 78.050 ;
        RECT 236.370 71.245 236.600 71.250 ;
        RECT 236.850 71.245 237.080 71.250 ;
        RECT 237.330 71.245 237.560 71.250 ;
        RECT 237.810 71.245 238.040 71.250 ;
        RECT 238.290 71.245 238.520 71.250 ;
        RECT 240.970 71.245 241.200 71.250 ;
        RECT 241.450 71.245 241.680 71.250 ;
        RECT 241.930 71.245 242.160 71.250 ;
        RECT 242.410 71.245 242.640 71.250 ;
        RECT 242.890 71.245 243.120 71.250 ;
        RECT 245.570 71.245 245.800 71.250 ;
        RECT 246.050 71.245 246.280 71.250 ;
        RECT 246.530 71.245 246.760 71.250 ;
        RECT 247.010 71.245 247.240 71.250 ;
        RECT 247.490 71.245 247.720 71.250 ;
        RECT 237.050 71.045 237.850 71.050 ;
        RECT 242.100 71.045 242.475 71.050 ;
        RECT 246.250 71.045 247.050 71.050 ;
        RECT 230.000 69.725 232.975 70.325 ;
        RECT 129.370 68.535 129.620 68.575 ;
        RECT 130.200 68.535 130.450 68.575 ;
        RECT 131.030 68.535 131.280 68.575 ;
        RECT 131.860 68.535 132.110 68.575 ;
        RECT 132.690 68.535 132.940 68.575 ;
        RECT 133.520 68.535 133.770 68.575 ;
        RECT 134.350 68.535 134.600 68.575 ;
        RECT 135.180 68.535 135.430 68.575 ;
        RECT 136.010 68.535 136.260 68.575 ;
        RECT 136.840 68.535 137.090 68.575 ;
        RECT 137.670 68.535 137.920 68.575 ;
        RECT 138.500 68.535 138.750 68.575 ;
        RECT 139.330 68.535 139.580 68.575 ;
        RECT 140.160 68.535 140.410 68.575 ;
        RECT 140.990 68.535 141.240 68.575 ;
        RECT 141.820 68.535 142.070 68.575 ;
        RECT 142.650 68.535 142.900 68.575 ;
        RECT 143.480 68.535 143.730 68.575 ;
        RECT 144.310 68.535 144.560 68.575 ;
        RECT 145.140 68.535 145.390 68.575 ;
        RECT 145.970 68.535 146.220 68.575 ;
        RECT 146.800 68.535 147.050 68.575 ;
        RECT 147.630 68.535 147.880 68.575 ;
        RECT 148.460 68.535 148.710 68.575 ;
        RECT 149.290 68.535 149.540 68.575 ;
        RECT 150.120 68.535 150.370 68.575 ;
        RECT 150.950 68.535 151.200 68.575 ;
        RECT 151.780 68.535 152.030 68.575 ;
        RECT 152.610 68.535 152.860 68.575 ;
        RECT 153.440 68.535 153.690 68.575 ;
        RECT 154.270 68.535 154.520 68.575 ;
        RECT 155.100 68.535 155.350 68.575 ;
        RECT 155.930 68.535 156.180 68.575 ;
        RECT 156.760 68.535 157.010 68.575 ;
        RECT 157.590 68.535 157.840 68.575 ;
        RECT 158.420 68.535 158.670 68.575 ;
        RECT 159.250 68.535 159.500 68.575 ;
        RECT 160.080 68.535 160.330 68.575 ;
        RECT 160.910 68.535 161.160 68.575 ;
        RECT 161.740 68.535 161.990 68.575 ;
        RECT 162.570 68.535 162.820 68.575 ;
        RECT 163.400 68.535 163.650 68.575 ;
        RECT 164.230 68.535 164.480 68.575 ;
        RECT 165.060 68.535 165.310 68.575 ;
        RECT 165.890 68.535 166.140 68.575 ;
        RECT 166.720 68.535 166.970 68.575 ;
        RECT 167.550 68.535 167.800 68.575 ;
        RECT 168.380 68.535 168.630 68.575 ;
        RECT 169.210 68.535 169.460 68.575 ;
        RECT 170.040 68.535 170.290 68.575 ;
        RECT 170.870 68.535 171.120 68.575 ;
        RECT 171.700 68.535 171.950 68.575 ;
        RECT 172.530 68.535 172.780 68.575 ;
        RECT 173.360 68.535 173.610 68.575 ;
        RECT 174.190 68.535 174.440 68.575 ;
        RECT 175.020 68.535 175.270 68.575 ;
        RECT 175.850 68.535 176.100 68.575 ;
        RECT 176.680 68.535 176.930 68.575 ;
        RECT 177.510 68.535 177.760 68.575 ;
        RECT 178.340 68.535 178.590 68.575 ;
        RECT 179.170 68.535 179.420 68.575 ;
        RECT 180.000 68.535 180.250 68.575 ;
        RECT 180.830 68.535 181.080 68.575 ;
        RECT 181.660 68.535 181.910 68.575 ;
        RECT 182.490 68.535 182.740 68.575 ;
        RECT 183.320 68.535 183.570 68.575 ;
        RECT 184.150 68.535 184.400 68.575 ;
        RECT 184.980 68.535 185.230 68.575 ;
        RECT 185.810 68.535 186.060 68.575 ;
        RECT 186.640 68.535 186.890 68.575 ;
        RECT 187.470 68.535 187.720 68.575 ;
        RECT 188.300 68.535 188.550 68.575 ;
        RECT 189.130 68.535 189.380 68.575 ;
        RECT 189.960 68.535 190.210 68.575 ;
        RECT 190.790 68.535 191.040 68.575 ;
        RECT 191.620 68.535 191.870 68.575 ;
        RECT 192.450 68.535 192.700 68.575 ;
        RECT 193.280 68.535 193.530 68.575 ;
        RECT 194.110 68.535 194.360 68.575 ;
        RECT 194.940 68.535 195.190 68.575 ;
        RECT 195.770 68.535 196.020 68.575 ;
        RECT 196.600 68.535 196.850 68.575 ;
        RECT 197.430 68.535 197.680 68.575 ;
        RECT 198.260 68.535 198.510 68.575 ;
        RECT 199.090 68.535 199.340 68.575 ;
        RECT 199.920 68.535 200.170 68.575 ;
        RECT 200.750 68.535 201.000 68.575 ;
        RECT 201.580 68.535 201.830 68.575 ;
        RECT 202.410 68.535 202.660 68.575 ;
        RECT 203.240 68.535 203.490 68.575 ;
        RECT 204.070 68.535 204.320 68.575 ;
        RECT 204.900 68.535 205.150 68.575 ;
        RECT 205.730 68.535 205.980 68.575 ;
        RECT 206.560 68.535 206.810 68.575 ;
        RECT 207.390 68.535 207.640 68.575 ;
        RECT 208.220 68.535 208.470 68.575 ;
        RECT 209.050 68.535 209.300 68.575 ;
        RECT 209.880 68.535 210.130 68.575 ;
        RECT 210.710 68.535 210.960 68.575 ;
        RECT 211.540 68.535 211.790 68.575 ;
        RECT 212.325 68.025 231.425 68.850 ;
        RECT 75.275 67.150 231.425 68.025 ;
        RECT 231.775 67.850 232.025 69.725 ;
        RECT 232.200 67.850 232.550 68.850 ;
        RECT 232.725 67.850 232.975 69.725 ;
        RECT 233.325 68.850 233.700 71.000 ;
        RECT 237.045 70.670 237.850 71.045 ;
        RECT 242.095 70.670 242.475 71.045 ;
        RECT 246.245 70.670 247.050 71.045 ;
        RECT 237.050 70.325 237.850 70.670 ;
        RECT 242.100 70.325 242.475 70.670 ;
        RECT 246.250 70.325 247.050 70.670 ;
        RECT 250.825 70.675 253.580 71.050 ;
        RECT 256.625 70.925 271.250 71.250 ;
        RECT 250.825 70.325 253.575 70.675 ;
        RECT 256.625 70.400 271.250 70.750 ;
        RECT 234.900 69.725 237.850 70.325 ;
        RECT 239.500 69.725 242.475 70.325 ;
        RECT 244.775 69.725 247.050 70.325 ;
        RECT 248.700 69.725 253.575 70.325 ;
        RECT 237.050 69.050 237.850 69.725 ;
        RECT 242.100 69.050 242.475 69.725 ;
        RECT 246.250 69.050 247.050 69.725 ;
        RECT 250.825 69.375 253.575 69.725 ;
        RECT 250.825 69.050 253.580 69.375 ;
        RECT 233.325 67.850 237.085 68.850 ;
        RECT 237.275 67.850 237.625 68.850 ;
        RECT 237.815 67.850 239.250 68.850 ;
        RECT 231.950 67.325 232.800 67.650 ;
        RECT 233.325 67.150 236.650 67.850 ;
        RECT 238.250 67.150 239.250 67.850 ;
        RECT 240.250 67.850 241.685 68.850 ;
        RECT 241.875 67.850 242.225 68.850 ;
        RECT 242.415 67.850 243.850 68.850 ;
        RECT 240.250 67.650 241.250 67.850 ;
        RECT 242.850 67.650 243.850 67.850 ;
        RECT 240.250 67.150 241.525 67.650 ;
        RECT 242.575 67.150 243.850 67.650 ;
        RECT 244.850 67.850 246.285 68.850 ;
        RECT 246.475 67.850 246.825 68.850 ;
        RECT 247.015 67.850 250.880 68.850 ;
        RECT 251.075 67.850 251.400 68.850 ;
        RECT 244.850 67.150 245.850 67.850 ;
        RECT 247.450 67.825 250.880 67.850 ;
        RECT 247.450 67.150 250.875 67.825 ;
        RECT 251.600 67.150 251.850 68.850 ;
        RECT 252.050 67.850 252.375 68.850 ;
        RECT 252.550 67.150 252.800 68.850 ;
        RECT 253.000 67.850 253.325 68.850 ;
        RECT 253.525 67.300 254.950 68.850 ;
        RECT 253.525 67.150 263.775 67.300 ;
        RECT 75.275 65.950 263.775 67.150 ;
        RECT 64.975 21.375 133.400 23.400 ;
        RECT 56.450 16.100 114.075 18.125 ;
        RECT 47.925 10.750 94.750 12.775 ;
        RECT 39.400 5.650 75.425 7.575 ;
      LAYER met2 ;
        RECT 56.450 215.100 127.600 217.150 ;
        RECT 56.450 137.250 58.475 215.100 ;
        RECT 138.275 213.850 139.100 214.450 ;
        RECT 135.525 210.575 136.350 211.175 ;
        RECT 132.775 207.300 133.600 207.900 ;
        RECT 130.000 204.050 130.825 204.650 ;
        RECT 75.275 156.550 81.175 158.225 ;
        RECT 111.925 151.275 113.050 201.100 ;
        RECT 127.675 157.325 128.825 157.375 ;
        RECT 180.125 157.325 181.250 201.100 ;
        RECT 127.675 155.250 181.250 157.325 ;
        RECT 179.900 151.250 180.350 153.375 ;
        RECT 180.650 151.250 181.250 155.250 ;
        RECT 216.400 158.500 266.400 159.850 ;
        RECT 212.800 151.300 214.125 153.325 ;
        RECT 216.400 150.600 223.825 158.500 ;
        RECT 232.675 154.650 233.025 157.900 ;
        RECT 237.275 154.650 237.625 157.900 ;
        RECT 239.425 154.975 240.075 157.825 ;
        RECT 241.875 154.675 242.225 157.900 ;
        RECT 244.025 154.975 244.675 157.825 ;
        RECT 232.675 154.300 233.625 154.650 ;
        RECT 237.275 154.300 238.225 154.650 ;
        RECT 241.875 154.300 242.825 154.675 ;
        RECT 246.475 154.650 246.825 157.900 ;
        RECT 246.475 154.300 247.425 154.650 ;
        RECT 233.025 153.975 233.625 154.300 ;
        RECT 237.625 153.975 238.225 154.300 ;
        RECT 242.225 153.975 242.825 154.300 ;
        RECT 246.825 153.975 247.425 154.300 ;
        RECT 251.075 153.975 251.400 157.900 ;
        RECT 252.050 153.975 252.375 157.900 ;
        RECT 253.000 153.975 253.325 157.900 ;
        RECT 233.025 153.375 235.400 153.975 ;
        RECT 237.625 153.375 240.000 153.975 ;
        RECT 241.175 153.375 241.975 153.975 ;
        RECT 242.225 153.375 243.925 153.975 ;
        RECT 245.775 153.375 246.575 153.975 ;
        RECT 246.825 153.375 249.200 153.975 ;
        RECT 251.075 153.375 256.000 153.975 ;
        RECT 233.025 153.075 233.625 153.375 ;
        RECT 237.625 153.075 238.225 153.375 ;
        RECT 242.225 153.075 242.825 153.375 ;
        RECT 246.825 153.075 247.425 153.375 ;
        RECT 232.675 152.725 233.625 153.075 ;
        RECT 237.275 152.725 238.225 153.075 ;
        RECT 232.675 151.500 233.025 152.725 ;
        RECT 75.025 149.900 226.125 150.600 ;
        RECT 234.825 150.525 235.475 152.425 ;
        RECT 237.275 151.500 237.625 152.725 ;
        RECT 241.875 152.700 242.825 153.075 ;
        RECT 246.475 152.725 247.425 153.075 ;
        RECT 241.875 151.500 242.225 152.700 ;
        RECT 246.475 151.500 246.825 152.725 ;
        RECT 248.625 150.525 249.275 152.425 ;
        RECT 251.075 151.500 251.400 153.375 ;
        RECT 252.050 151.500 252.375 153.375 ;
        RECT 253.000 151.500 253.325 153.375 ;
        RECT 255.400 153.000 256.000 153.375 ;
        RECT 255.400 152.400 271.250 153.000 ;
        RECT 257.300 150.950 259.050 152.125 ;
        RECT 259.700 150.950 270.575 152.125 ;
        RECT 65.000 149.150 226.125 149.900 ;
        RECT 242.450 149.750 246.825 150.400 ;
        RECT 65.000 148.175 75.050 149.150 ;
        RECT 231.950 148.800 233.700 149.175 ;
        RECT 84.330 147.920 225.105 148.670 ;
        RECT 78.305 137.620 79.105 146.820 ;
        RECT 80.855 137.620 81.655 146.820 ;
        RECT 84.330 137.620 85.080 147.920 ;
        RECT 56.450 136.000 73.525 137.250 ;
        RECT 78.305 135.620 85.080 137.620 ;
        RECT 85.680 135.845 86.655 137.395 ;
        RECT 78.305 132.470 79.105 135.620 ;
        RECT 80.855 132.470 81.655 135.620 ;
        RECT 87.030 131.420 87.880 146.820 ;
        RECT 89.055 137.620 89.855 146.820 ;
        RECT 91.630 137.620 92.430 146.820 ;
        RECT 94.205 137.620 95.005 146.820 ;
        RECT 96.855 141.820 99.355 143.370 ;
        RECT 96.855 137.620 98.405 141.820 ;
        RECT 89.055 135.620 98.405 137.620 ;
        RECT 99.005 135.845 99.980 137.395 ;
        RECT 89.055 132.470 89.855 135.620 ;
        RECT 91.630 132.470 92.430 135.620 ;
        RECT 94.205 132.470 95.005 135.620 ;
        RECT 100.355 131.420 101.205 146.820 ;
        RECT 102.380 137.620 103.180 146.820 ;
        RECT 104.955 137.620 105.755 146.820 ;
        RECT 107.530 137.620 108.330 146.820 ;
        RECT 110.180 141.820 112.680 143.370 ;
        RECT 110.180 137.620 111.730 141.820 ;
        RECT 102.380 137.395 111.730 137.620 ;
        RECT 102.380 135.845 113.305 137.395 ;
        RECT 102.380 135.620 111.730 135.845 ;
        RECT 102.380 132.470 103.180 135.620 ;
        RECT 104.955 132.470 105.755 135.620 ;
        RECT 107.530 132.470 108.330 135.620 ;
        RECT 113.680 131.420 114.530 146.820 ;
        RECT 115.705 137.620 116.505 146.820 ;
        RECT 118.255 137.620 119.055 146.820 ;
        RECT 115.705 135.620 122.455 137.620 ;
        RECT 123.080 135.845 124.055 137.395 ;
        RECT 115.705 132.470 116.505 135.620 ;
        RECT 118.255 132.470 119.055 135.620 ;
        RECT 120.905 134.645 122.455 135.620 ;
        RECT 120.905 133.095 123.430 134.645 ;
        RECT 124.430 131.420 125.280 146.820 ;
        RECT 126.455 137.620 127.255 146.820 ;
        RECT 129.030 137.620 129.830 146.820 ;
        RECT 131.605 137.620 132.405 146.820 ;
        RECT 134.230 141.820 136.755 143.370 ;
        RECT 134.230 137.620 135.780 141.820 ;
        RECT 126.455 135.620 135.780 137.620 ;
        RECT 136.405 135.845 137.380 137.395 ;
        RECT 126.455 132.470 127.255 135.620 ;
        RECT 129.030 132.470 129.830 135.620 ;
        RECT 131.605 132.470 132.405 135.620 ;
        RECT 137.755 131.420 138.605 146.820 ;
        RECT 139.780 137.620 140.580 146.820 ;
        RECT 142.355 137.620 143.155 146.820 ;
        RECT 144.930 137.620 145.730 146.820 ;
        RECT 139.780 135.620 149.105 137.620 ;
        RECT 149.730 135.845 150.705 137.395 ;
        RECT 139.780 132.470 140.580 135.620 ;
        RECT 142.355 132.470 143.155 135.620 ;
        RECT 144.930 132.470 145.730 135.620 ;
        RECT 147.555 134.645 149.105 135.620 ;
        RECT 147.555 133.095 150.080 134.645 ;
        RECT 151.080 131.420 151.930 146.820 ;
        RECT 153.105 137.620 153.905 146.820 ;
        RECT 155.680 137.620 156.480 146.820 ;
        RECT 158.255 137.620 159.055 146.820 ;
        RECT 160.880 141.820 163.405 143.370 ;
        RECT 160.880 137.620 162.430 141.820 ;
        RECT 153.105 135.620 162.430 137.620 ;
        RECT 163.055 135.845 164.030 137.395 ;
        RECT 153.105 132.470 153.905 135.620 ;
        RECT 155.680 132.470 156.480 135.620 ;
        RECT 158.255 132.470 159.055 135.620 ;
        RECT 164.405 131.420 165.255 146.820 ;
        RECT 166.430 137.620 167.230 146.820 ;
        RECT 169.005 137.620 169.805 146.820 ;
        RECT 171.580 137.620 172.380 146.820 ;
        RECT 166.430 135.620 175.755 137.620 ;
        RECT 176.380 135.845 177.355 137.395 ;
        RECT 166.430 132.470 167.230 135.620 ;
        RECT 169.005 132.470 169.805 135.620 ;
        RECT 171.580 132.470 172.380 135.620 ;
        RECT 177.730 131.420 178.580 146.820 ;
        RECT 179.755 137.620 180.555 146.820 ;
        RECT 182.330 137.620 183.130 146.820 ;
        RECT 184.905 137.620 185.705 146.820 ;
        RECT 187.530 138.270 190.055 139.820 ;
        RECT 187.530 137.620 189.080 138.270 ;
        RECT 179.755 135.620 189.080 137.620 ;
        RECT 189.705 135.845 190.680 137.395 ;
        RECT 179.755 132.470 180.555 135.620 ;
        RECT 182.330 132.470 183.130 135.620 ;
        RECT 184.905 132.470 185.705 135.620 ;
        RECT 191.055 131.420 191.905 146.820 ;
        RECT 193.080 137.620 193.880 146.820 ;
        RECT 195.630 137.620 196.430 146.820 ;
        RECT 193.080 135.620 199.555 137.620 ;
        RECT 200.455 135.845 201.430 137.395 ;
        RECT 193.080 132.470 193.880 135.620 ;
        RECT 195.630 132.470 196.430 135.620 ;
        RECT 201.805 131.420 202.655 146.820 ;
        RECT 203.830 137.620 204.630 146.820 ;
        RECT 206.405 137.620 207.205 146.820 ;
        RECT 208.980 137.620 209.780 146.820 ;
        RECT 211.605 141.820 214.130 143.370 ;
        RECT 211.605 137.620 213.155 141.820 ;
        RECT 203.830 135.620 213.155 137.620 ;
        RECT 213.780 135.845 214.755 137.395 ;
        RECT 203.830 132.470 204.630 135.620 ;
        RECT 206.405 132.470 207.205 135.620 ;
        RECT 208.980 132.470 209.780 135.620 ;
        RECT 215.130 131.420 215.980 146.820 ;
        RECT 217.155 137.620 217.955 146.820 ;
        RECT 219.730 137.620 220.530 146.820 ;
        RECT 222.305 137.620 223.105 146.820 ;
        RECT 224.880 141.820 227.455 143.370 ;
        RECT 224.880 137.620 226.430 141.820 ;
        RECT 228.675 139.800 229.275 144.250 ;
        RECT 231.050 142.025 231.425 148.625 ;
        RECT 232.200 144.675 232.550 148.625 ;
        RECT 233.325 144.925 233.700 148.800 ;
        RECT 237.275 145.350 237.625 148.600 ;
        RECT 239.425 145.675 240.075 148.525 ;
        RECT 241.875 145.375 242.225 148.600 ;
        RECT 244.025 145.675 244.675 148.525 ;
        RECT 237.275 145.000 238.225 145.350 ;
        RECT 241.875 145.000 242.825 145.375 ;
        RECT 246.475 145.350 246.825 148.600 ;
        RECT 246.475 145.000 247.425 145.350 ;
        RECT 237.625 144.675 238.225 145.000 ;
        RECT 242.225 144.675 242.825 145.000 ;
        RECT 246.825 144.675 247.425 145.000 ;
        RECT 251.075 144.675 251.400 148.600 ;
        RECT 252.050 144.675 252.375 148.600 ;
        RECT 253.000 144.675 253.325 148.600 ;
        RECT 255.400 147.675 258.700 148.325 ;
        RECT 255.400 144.675 256.000 147.675 ;
        RECT 259.200 146.450 268.225 150.325 ;
        RECT 257.300 145.750 259.025 146.150 ;
        RECT 259.700 145.750 270.575 146.150 ;
        RECT 232.200 144.075 235.400 144.675 ;
        RECT 237.625 144.075 240.000 144.675 ;
        RECT 241.175 144.075 241.975 144.675 ;
        RECT 242.225 144.075 243.925 144.675 ;
        RECT 245.775 144.075 246.575 144.675 ;
        RECT 246.825 144.075 249.200 144.675 ;
        RECT 251.075 144.075 256.000 144.675 ;
        RECT 232.200 142.200 232.550 144.075 ;
        RECT 237.625 143.775 238.225 144.075 ;
        RECT 242.225 143.775 242.825 144.075 ;
        RECT 246.825 143.775 247.425 144.075 ;
        RECT 237.275 143.425 238.225 143.775 ;
        RECT 231.050 141.650 232.800 142.025 ;
        RECT 234.825 141.225 235.475 143.125 ;
        RECT 237.275 142.200 237.625 143.425 ;
        RECT 241.875 143.400 242.825 143.775 ;
        RECT 246.475 143.425 247.425 143.775 ;
        RECT 241.875 142.200 242.225 143.400 ;
        RECT 246.475 142.200 246.825 143.425 ;
        RECT 248.625 141.225 249.275 143.125 ;
        RECT 251.075 142.200 251.400 144.075 ;
        RECT 252.050 142.200 252.375 144.075 ;
        RECT 253.000 142.200 253.325 144.075 ;
        RECT 258.350 140.300 261.450 141.650 ;
        RECT 228.675 139.200 230.600 139.800 ;
        RECT 263.300 137.650 266.400 139.000 ;
        RECT 217.155 135.620 226.430 137.620 ;
        RECT 217.155 132.470 217.955 135.620 ;
        RECT 219.730 132.470 220.530 135.620 ;
        RECT 222.305 132.470 223.105 135.620 ;
        RECT 232.675 133.800 233.025 137.050 ;
        RECT 237.275 133.800 237.625 137.050 ;
        RECT 239.425 134.125 240.075 136.975 ;
        RECT 241.875 133.825 242.225 137.050 ;
        RECT 244.025 134.125 244.675 136.975 ;
        RECT 232.675 133.450 233.625 133.800 ;
        RECT 237.275 133.450 238.225 133.800 ;
        RECT 241.875 133.450 242.825 133.825 ;
        RECT 246.475 133.800 246.825 137.050 ;
        RECT 246.475 133.450 247.425 133.800 ;
        RECT 233.025 133.125 233.625 133.450 ;
        RECT 237.625 133.125 238.225 133.450 ;
        RECT 242.225 133.125 242.825 133.450 ;
        RECT 246.825 133.125 247.425 133.450 ;
        RECT 251.075 133.125 251.400 137.050 ;
        RECT 252.050 133.125 252.375 137.050 ;
        RECT 253.000 133.125 253.325 137.050 ;
        RECT 233.025 132.525 235.400 133.125 ;
        RECT 237.625 132.525 240.000 133.125 ;
        RECT 241.175 132.525 241.975 133.125 ;
        RECT 242.225 132.525 243.925 133.125 ;
        RECT 245.775 132.525 246.575 133.125 ;
        RECT 246.825 132.525 249.200 133.125 ;
        RECT 251.075 132.525 256.000 133.125 ;
        RECT 233.025 132.225 233.625 132.525 ;
        RECT 237.625 132.225 238.225 132.525 ;
        RECT 242.225 132.225 242.825 132.525 ;
        RECT 246.825 132.225 247.425 132.525 ;
        RECT 232.675 131.875 233.625 132.225 ;
        RECT 237.275 131.875 238.225 132.225 ;
        RECT 75.275 129.450 81.175 131.125 ;
        RECT 87.030 130.670 97.005 131.420 ;
        RECT 100.355 130.670 110.330 131.420 ;
        RECT 113.680 130.670 121.030 131.420 ;
        RECT 124.430 130.670 134.405 131.420 ;
        RECT 137.755 130.670 147.730 131.420 ;
        RECT 151.080 130.670 161.055 131.420 ;
        RECT 164.405 130.670 174.380 131.420 ;
        RECT 177.730 130.670 187.705 131.420 ;
        RECT 191.055 130.670 198.405 131.420 ;
        RECT 201.805 130.670 211.780 131.420 ;
        RECT 215.130 130.670 225.105 131.420 ;
        RECT 232.675 130.650 233.025 131.875 ;
        RECT 234.825 129.675 235.475 131.575 ;
        RECT 237.275 130.650 237.625 131.875 ;
        RECT 241.875 131.850 242.825 132.225 ;
        RECT 246.475 131.875 247.425 132.225 ;
        RECT 241.875 130.650 242.225 131.850 ;
        RECT 246.475 130.650 246.825 131.875 ;
        RECT 248.625 129.675 249.275 131.575 ;
        RECT 251.075 130.650 251.400 132.525 ;
        RECT 252.050 130.650 252.375 132.525 ;
        RECT 253.000 130.650 253.325 132.525 ;
        RECT 255.400 132.150 256.000 132.525 ;
        RECT 255.400 131.550 271.250 132.150 ;
        RECT 257.300 130.100 259.050 131.275 ;
        RECT 259.700 130.100 270.575 131.275 ;
        RECT 242.450 128.900 246.825 129.550 ;
        RECT 111.925 126.075 113.050 127.200 ;
        RECT 179.900 126.025 180.350 128.150 ;
        RECT 180.650 124.150 181.250 128.150 ;
        RECT 212.800 126.075 214.125 128.100 ;
        RECT 231.950 127.950 233.700 128.325 ;
        RECT 75.275 121.175 81.175 122.850 ;
        RECT 127.675 122.025 207.800 124.150 ;
        RECT 231.050 121.175 231.425 127.775 ;
        RECT 232.200 123.825 232.550 127.775 ;
        RECT 233.325 124.075 233.700 127.950 ;
        RECT 237.275 124.500 237.625 127.750 ;
        RECT 239.425 124.825 240.075 127.675 ;
        RECT 241.875 124.525 242.225 127.750 ;
        RECT 244.025 124.825 244.675 127.675 ;
        RECT 237.275 124.150 238.225 124.500 ;
        RECT 241.875 124.150 242.825 124.525 ;
        RECT 246.475 124.500 246.825 127.750 ;
        RECT 246.475 124.150 247.425 124.500 ;
        RECT 237.625 123.825 238.225 124.150 ;
        RECT 242.225 123.825 242.825 124.150 ;
        RECT 246.825 123.825 247.425 124.150 ;
        RECT 251.075 123.825 251.400 127.750 ;
        RECT 252.050 123.825 252.375 127.750 ;
        RECT 253.000 123.825 253.325 127.750 ;
        RECT 255.125 126.800 258.425 127.450 ;
        RECT 255.125 123.825 255.725 126.800 ;
        RECT 259.200 125.600 268.225 129.475 ;
        RECT 257.300 124.900 259.025 125.300 ;
        RECT 259.700 124.900 270.575 125.300 ;
        RECT 232.200 123.225 235.400 123.825 ;
        RECT 237.625 123.225 240.000 123.825 ;
        RECT 241.175 123.225 241.975 123.825 ;
        RECT 242.225 123.225 243.925 123.825 ;
        RECT 245.775 123.225 246.575 123.825 ;
        RECT 246.825 123.225 249.200 123.825 ;
        RECT 251.075 123.225 256.000 123.825 ;
        RECT 232.200 121.350 232.550 123.225 ;
        RECT 237.625 122.925 238.225 123.225 ;
        RECT 242.225 122.925 242.825 123.225 ;
        RECT 246.825 122.925 247.425 123.225 ;
        RECT 237.275 122.575 238.225 122.925 ;
        RECT 231.050 120.800 232.800 121.175 ;
        RECT 234.825 120.375 235.475 122.275 ;
        RECT 237.275 121.350 237.625 122.575 ;
        RECT 241.875 122.550 242.825 122.925 ;
        RECT 246.475 122.575 247.425 122.925 ;
        RECT 241.875 121.350 242.225 122.550 ;
        RECT 246.475 121.350 246.825 122.575 ;
        RECT 248.625 120.375 249.275 122.275 ;
        RECT 251.075 121.350 251.400 123.225 ;
        RECT 252.050 121.350 252.375 123.225 ;
        RECT 253.000 121.350 253.325 123.225 ;
        RECT 260.675 119.450 263.775 120.800 ;
        RECT 75.275 110.200 81.175 111.300 ;
        RECT 56.450 104.275 81.175 110.200 ;
        RECT 75.275 103.050 81.175 104.275 ;
        RECT 216.400 105.000 266.400 106.350 ;
        RECT 127.675 103.825 128.825 103.875 ;
        RECT 127.675 101.750 207.800 103.825 ;
        RECT 111.925 98.775 113.050 99.825 ;
        RECT 179.900 97.750 180.350 99.875 ;
        RECT 180.650 97.750 181.250 101.750 ;
        RECT 212.800 97.800 214.125 99.825 ;
        RECT 216.400 97.100 223.825 105.000 ;
        RECT 232.675 101.150 233.025 104.400 ;
        RECT 237.275 101.150 237.625 104.400 ;
        RECT 239.425 101.475 240.075 104.325 ;
        RECT 241.875 101.175 242.225 104.400 ;
        RECT 244.025 101.475 244.675 104.325 ;
        RECT 232.675 100.800 233.625 101.150 ;
        RECT 237.275 100.800 238.225 101.150 ;
        RECT 241.875 100.800 242.825 101.175 ;
        RECT 246.475 101.150 246.825 104.400 ;
        RECT 246.475 100.800 247.425 101.150 ;
        RECT 233.025 100.475 233.625 100.800 ;
        RECT 237.625 100.475 238.225 100.800 ;
        RECT 242.225 100.475 242.825 100.800 ;
        RECT 246.825 100.475 247.425 100.800 ;
        RECT 251.075 100.475 251.400 104.400 ;
        RECT 252.050 100.475 252.375 104.400 ;
        RECT 253.000 100.475 253.325 104.400 ;
        RECT 233.025 99.875 235.400 100.475 ;
        RECT 237.625 99.875 240.000 100.475 ;
        RECT 241.175 99.875 241.975 100.475 ;
        RECT 242.225 99.875 243.925 100.475 ;
        RECT 245.775 99.875 246.575 100.475 ;
        RECT 246.825 99.875 249.200 100.475 ;
        RECT 251.075 99.875 256.000 100.475 ;
        RECT 233.025 99.575 233.625 99.875 ;
        RECT 237.625 99.575 238.225 99.875 ;
        RECT 242.225 99.575 242.825 99.875 ;
        RECT 246.825 99.575 247.425 99.875 ;
        RECT 232.675 99.225 233.625 99.575 ;
        RECT 237.275 99.225 238.225 99.575 ;
        RECT 232.675 98.000 233.025 99.225 ;
        RECT 75.025 96.400 226.125 97.100 ;
        RECT 234.825 97.025 235.475 98.925 ;
        RECT 237.275 98.000 237.625 99.225 ;
        RECT 241.875 99.200 242.825 99.575 ;
        RECT 246.475 99.225 247.425 99.575 ;
        RECT 241.875 98.000 242.225 99.200 ;
        RECT 246.475 98.000 246.825 99.225 ;
        RECT 248.625 97.025 249.275 98.925 ;
        RECT 251.075 98.000 251.400 99.875 ;
        RECT 252.050 98.000 252.375 99.875 ;
        RECT 253.000 98.000 253.325 99.875 ;
        RECT 255.400 99.500 256.000 99.875 ;
        RECT 255.400 98.900 271.250 99.500 ;
        RECT 257.300 97.450 259.050 98.625 ;
        RECT 259.700 97.450 270.575 98.625 ;
        RECT 65.000 95.650 226.125 96.400 ;
        RECT 242.450 96.250 246.825 96.900 ;
        RECT 65.000 94.675 75.050 95.650 ;
        RECT 231.950 95.300 233.700 95.675 ;
        RECT 84.330 94.420 225.105 95.170 ;
        RECT 78.305 84.120 79.105 93.320 ;
        RECT 80.855 84.120 81.655 93.320 ;
        RECT 84.330 84.120 85.080 94.420 ;
        RECT 72.650 82.500 73.525 83.750 ;
        RECT 78.305 82.120 85.080 84.120 ;
        RECT 85.680 82.345 86.655 83.895 ;
        RECT 78.305 78.970 79.105 82.120 ;
        RECT 80.855 78.970 81.655 82.120 ;
        RECT 87.030 77.920 87.880 93.320 ;
        RECT 89.055 84.120 89.855 93.320 ;
        RECT 91.630 84.120 92.430 93.320 ;
        RECT 94.205 84.120 95.005 93.320 ;
        RECT 96.855 88.320 99.355 89.870 ;
        RECT 96.855 84.120 98.405 88.320 ;
        RECT 89.055 82.120 98.405 84.120 ;
        RECT 99.005 82.345 99.980 83.895 ;
        RECT 89.055 78.970 89.855 82.120 ;
        RECT 91.630 78.970 92.430 82.120 ;
        RECT 94.205 78.970 95.005 82.120 ;
        RECT 100.355 77.920 101.205 93.320 ;
        RECT 102.380 84.120 103.180 93.320 ;
        RECT 104.955 84.120 105.755 93.320 ;
        RECT 107.530 84.120 108.330 93.320 ;
        RECT 110.180 88.320 112.680 89.870 ;
        RECT 110.180 84.120 111.730 88.320 ;
        RECT 102.380 83.895 111.730 84.120 ;
        RECT 102.380 82.345 113.305 83.895 ;
        RECT 102.380 82.120 111.730 82.345 ;
        RECT 102.380 78.970 103.180 82.120 ;
        RECT 104.955 78.970 105.755 82.120 ;
        RECT 107.530 78.970 108.330 82.120 ;
        RECT 113.680 77.920 114.530 93.320 ;
        RECT 115.705 84.120 116.505 93.320 ;
        RECT 118.255 84.120 119.055 93.320 ;
        RECT 115.705 82.120 122.455 84.120 ;
        RECT 123.080 82.345 124.055 83.895 ;
        RECT 115.705 78.970 116.505 82.120 ;
        RECT 118.255 78.970 119.055 82.120 ;
        RECT 120.905 81.145 122.455 82.120 ;
        RECT 120.905 79.595 123.430 81.145 ;
        RECT 124.430 77.920 125.280 93.320 ;
        RECT 126.455 84.120 127.255 93.320 ;
        RECT 129.030 84.120 129.830 93.320 ;
        RECT 131.605 84.120 132.405 93.320 ;
        RECT 134.230 88.320 136.755 89.870 ;
        RECT 134.230 84.120 135.780 88.320 ;
        RECT 126.455 82.120 135.780 84.120 ;
        RECT 136.405 82.345 137.380 83.895 ;
        RECT 126.455 78.970 127.255 82.120 ;
        RECT 129.030 78.970 129.830 82.120 ;
        RECT 131.605 78.970 132.405 82.120 ;
        RECT 137.755 77.920 138.605 93.320 ;
        RECT 139.780 84.120 140.580 93.320 ;
        RECT 142.355 84.120 143.155 93.320 ;
        RECT 144.930 84.120 145.730 93.320 ;
        RECT 139.780 82.120 149.105 84.120 ;
        RECT 149.730 82.345 150.705 83.895 ;
        RECT 139.780 78.970 140.580 82.120 ;
        RECT 142.355 78.970 143.155 82.120 ;
        RECT 144.930 78.970 145.730 82.120 ;
        RECT 147.555 81.145 149.105 82.120 ;
        RECT 147.555 79.595 150.080 81.145 ;
        RECT 151.080 77.920 151.930 93.320 ;
        RECT 153.105 84.120 153.905 93.320 ;
        RECT 155.680 84.120 156.480 93.320 ;
        RECT 158.255 84.120 159.055 93.320 ;
        RECT 160.880 88.320 163.405 89.870 ;
        RECT 160.880 84.120 162.430 88.320 ;
        RECT 153.105 82.120 162.430 84.120 ;
        RECT 163.055 82.345 164.030 83.895 ;
        RECT 153.105 78.970 153.905 82.120 ;
        RECT 155.680 78.970 156.480 82.120 ;
        RECT 158.255 78.970 159.055 82.120 ;
        RECT 164.405 77.920 165.255 93.320 ;
        RECT 166.430 84.120 167.230 93.320 ;
        RECT 169.005 84.120 169.805 93.320 ;
        RECT 171.580 84.120 172.380 93.320 ;
        RECT 166.430 82.120 175.755 84.120 ;
        RECT 176.380 82.345 177.355 83.895 ;
        RECT 166.430 78.970 167.230 82.120 ;
        RECT 169.005 78.970 169.805 82.120 ;
        RECT 171.580 78.970 172.380 82.120 ;
        RECT 177.730 77.920 178.580 93.320 ;
        RECT 179.755 84.120 180.555 93.320 ;
        RECT 182.330 84.120 183.130 93.320 ;
        RECT 184.905 84.120 185.705 93.320 ;
        RECT 187.530 84.770 190.055 86.320 ;
        RECT 187.530 84.120 189.080 84.770 ;
        RECT 179.755 82.120 189.080 84.120 ;
        RECT 189.705 82.345 190.680 83.895 ;
        RECT 179.755 78.970 180.555 82.120 ;
        RECT 182.330 78.970 183.130 82.120 ;
        RECT 184.905 78.970 185.705 82.120 ;
        RECT 191.055 77.920 191.905 93.320 ;
        RECT 193.080 84.120 193.880 93.320 ;
        RECT 195.630 84.120 196.430 93.320 ;
        RECT 193.080 82.120 199.555 84.120 ;
        RECT 200.455 82.345 201.430 83.895 ;
        RECT 193.080 78.970 193.880 82.120 ;
        RECT 195.630 78.970 196.430 82.120 ;
        RECT 201.805 77.920 202.655 93.320 ;
        RECT 203.830 84.120 204.630 93.320 ;
        RECT 206.405 84.120 207.205 93.320 ;
        RECT 208.980 84.120 209.780 93.320 ;
        RECT 211.605 88.320 214.130 89.870 ;
        RECT 211.605 84.120 213.155 88.320 ;
        RECT 203.830 82.120 213.155 84.120 ;
        RECT 213.780 82.345 214.755 83.895 ;
        RECT 203.830 78.970 204.630 82.120 ;
        RECT 206.405 78.970 207.205 82.120 ;
        RECT 208.980 78.970 209.780 82.120 ;
        RECT 215.130 77.920 215.980 93.320 ;
        RECT 217.155 84.120 217.955 93.320 ;
        RECT 219.730 84.120 220.530 93.320 ;
        RECT 222.305 84.120 223.105 93.320 ;
        RECT 224.880 88.320 227.455 89.870 ;
        RECT 224.880 84.120 226.430 88.320 ;
        RECT 228.675 86.300 229.275 90.750 ;
        RECT 231.050 88.525 231.425 95.125 ;
        RECT 232.200 91.175 232.550 95.125 ;
        RECT 233.325 91.425 233.700 95.300 ;
        RECT 237.275 91.850 237.625 95.100 ;
        RECT 239.425 92.175 240.075 95.025 ;
        RECT 241.875 91.875 242.225 95.100 ;
        RECT 244.025 92.175 244.675 95.025 ;
        RECT 237.275 91.500 238.225 91.850 ;
        RECT 241.875 91.500 242.825 91.875 ;
        RECT 246.475 91.850 246.825 95.100 ;
        RECT 246.475 91.500 247.425 91.850 ;
        RECT 237.625 91.175 238.225 91.500 ;
        RECT 242.225 91.175 242.825 91.500 ;
        RECT 246.825 91.175 247.425 91.500 ;
        RECT 251.075 91.175 251.400 95.100 ;
        RECT 252.050 91.175 252.375 95.100 ;
        RECT 253.000 91.175 253.325 95.100 ;
        RECT 255.400 94.175 258.700 94.825 ;
        RECT 255.400 91.175 256.000 94.175 ;
        RECT 259.200 92.950 268.225 96.825 ;
        RECT 257.300 92.250 259.025 92.650 ;
        RECT 259.700 92.250 270.575 92.650 ;
        RECT 232.200 90.575 235.400 91.175 ;
        RECT 237.625 90.575 240.000 91.175 ;
        RECT 241.175 90.575 241.975 91.175 ;
        RECT 242.225 90.575 243.925 91.175 ;
        RECT 245.775 90.575 246.575 91.175 ;
        RECT 246.825 90.575 249.200 91.175 ;
        RECT 251.075 90.575 256.000 91.175 ;
        RECT 232.200 88.700 232.550 90.575 ;
        RECT 237.625 90.275 238.225 90.575 ;
        RECT 242.225 90.275 242.825 90.575 ;
        RECT 246.825 90.275 247.425 90.575 ;
        RECT 237.275 89.925 238.225 90.275 ;
        RECT 231.050 88.150 232.800 88.525 ;
        RECT 234.825 87.725 235.475 89.625 ;
        RECT 237.275 88.700 237.625 89.925 ;
        RECT 241.875 89.900 242.825 90.275 ;
        RECT 246.475 89.925 247.425 90.275 ;
        RECT 241.875 88.700 242.225 89.900 ;
        RECT 246.475 88.700 246.825 89.925 ;
        RECT 248.625 87.725 249.275 89.625 ;
        RECT 251.075 88.700 251.400 90.575 ;
        RECT 252.050 88.700 252.375 90.575 ;
        RECT 253.000 88.700 253.325 90.575 ;
        RECT 258.350 86.800 261.450 88.150 ;
        RECT 228.675 85.700 230.600 86.300 ;
        RECT 263.300 84.150 266.400 85.500 ;
        RECT 217.155 82.120 226.430 84.120 ;
        RECT 217.155 78.970 217.955 82.120 ;
        RECT 219.730 78.970 220.530 82.120 ;
        RECT 222.305 78.970 223.105 82.120 ;
        RECT 232.675 80.300 233.025 83.550 ;
        RECT 237.275 80.300 237.625 83.550 ;
        RECT 239.425 80.625 240.075 83.475 ;
        RECT 241.875 80.325 242.225 83.550 ;
        RECT 244.025 80.625 244.675 83.475 ;
        RECT 232.675 79.950 233.625 80.300 ;
        RECT 237.275 79.950 238.225 80.300 ;
        RECT 241.875 79.950 242.825 80.325 ;
        RECT 246.475 80.300 246.825 83.550 ;
        RECT 246.475 79.950 247.425 80.300 ;
        RECT 233.025 79.625 233.625 79.950 ;
        RECT 237.625 79.625 238.225 79.950 ;
        RECT 242.225 79.625 242.825 79.950 ;
        RECT 246.825 79.625 247.425 79.950 ;
        RECT 251.075 79.625 251.400 83.550 ;
        RECT 252.050 79.625 252.375 83.550 ;
        RECT 253.000 79.625 253.325 83.550 ;
        RECT 233.025 79.025 235.400 79.625 ;
        RECT 237.625 79.025 240.000 79.625 ;
        RECT 241.175 79.025 241.975 79.625 ;
        RECT 242.225 79.025 243.925 79.625 ;
        RECT 245.775 79.025 246.575 79.625 ;
        RECT 246.825 79.025 249.200 79.625 ;
        RECT 251.075 79.025 256.000 79.625 ;
        RECT 233.025 78.725 233.625 79.025 ;
        RECT 237.625 78.725 238.225 79.025 ;
        RECT 242.225 78.725 242.825 79.025 ;
        RECT 246.825 78.725 247.425 79.025 ;
        RECT 232.675 78.375 233.625 78.725 ;
        RECT 237.275 78.375 238.225 78.725 ;
        RECT 75.275 75.950 81.175 77.625 ;
        RECT 87.030 77.170 97.005 77.920 ;
        RECT 100.355 77.170 110.330 77.920 ;
        RECT 113.680 77.170 121.030 77.920 ;
        RECT 124.430 77.170 134.405 77.920 ;
        RECT 137.755 77.170 147.730 77.920 ;
        RECT 151.080 77.170 161.055 77.920 ;
        RECT 164.405 77.170 174.380 77.920 ;
        RECT 177.730 77.170 187.705 77.920 ;
        RECT 191.055 77.170 198.405 77.920 ;
        RECT 201.805 77.170 211.780 77.920 ;
        RECT 215.130 77.170 225.105 77.920 ;
        RECT 232.675 77.150 233.025 78.375 ;
        RECT 234.825 76.175 235.475 78.075 ;
        RECT 237.275 77.150 237.625 78.375 ;
        RECT 241.875 78.350 242.825 78.725 ;
        RECT 246.475 78.375 247.425 78.725 ;
        RECT 241.875 77.150 242.225 78.350 ;
        RECT 246.475 77.150 246.825 78.375 ;
        RECT 248.625 76.175 249.275 78.075 ;
        RECT 251.075 77.150 251.400 79.025 ;
        RECT 252.050 77.150 252.375 79.025 ;
        RECT 253.000 77.150 253.325 79.025 ;
        RECT 255.400 78.650 256.000 79.025 ;
        RECT 255.400 78.050 271.250 78.650 ;
        RECT 257.300 76.600 259.050 77.775 ;
        RECT 259.700 76.600 270.575 77.775 ;
        RECT 242.450 75.400 246.825 76.050 ;
        RECT 75.275 67.675 81.175 69.350 ;
        RECT 111.925 25.000 113.050 74.625 ;
        RECT 179.900 72.525 180.350 74.650 ;
        RECT 180.650 70.650 181.250 74.650 ;
        RECT 212.800 72.575 214.125 74.600 ;
        RECT 231.950 74.450 233.700 74.825 ;
        RECT 127.675 68.525 181.250 70.650 ;
        RECT 180.125 25.000 181.250 68.525 ;
        RECT 231.050 67.675 231.425 74.275 ;
        RECT 232.200 70.325 232.550 74.275 ;
        RECT 233.325 70.575 233.700 74.450 ;
        RECT 237.275 71.000 237.625 74.250 ;
        RECT 239.425 71.325 240.075 74.175 ;
        RECT 241.875 71.025 242.225 74.250 ;
        RECT 244.025 71.325 244.675 74.175 ;
        RECT 237.275 70.650 238.225 71.000 ;
        RECT 241.875 70.650 242.825 71.025 ;
        RECT 246.475 71.000 246.825 74.250 ;
        RECT 246.475 70.650 247.425 71.000 ;
        RECT 237.625 70.325 238.225 70.650 ;
        RECT 242.225 70.325 242.825 70.650 ;
        RECT 246.825 70.325 247.425 70.650 ;
        RECT 251.075 70.325 251.400 74.250 ;
        RECT 252.050 70.325 252.375 74.250 ;
        RECT 253.000 70.325 253.325 74.250 ;
        RECT 255.125 73.300 258.425 73.950 ;
        RECT 255.125 70.325 255.725 73.300 ;
        RECT 259.200 72.100 268.225 75.975 ;
        RECT 257.300 71.400 259.025 71.800 ;
        RECT 259.700 71.400 270.575 71.800 ;
        RECT 232.200 69.725 235.400 70.325 ;
        RECT 237.625 69.725 240.000 70.325 ;
        RECT 241.175 69.725 241.975 70.325 ;
        RECT 242.225 69.725 243.925 70.325 ;
        RECT 245.775 69.725 246.575 70.325 ;
        RECT 246.825 69.725 249.200 70.325 ;
        RECT 251.075 69.725 256.000 70.325 ;
        RECT 232.200 67.850 232.550 69.725 ;
        RECT 237.625 69.425 238.225 69.725 ;
        RECT 242.225 69.425 242.825 69.725 ;
        RECT 246.825 69.425 247.425 69.725 ;
        RECT 237.275 69.075 238.225 69.425 ;
        RECT 231.050 67.300 232.800 67.675 ;
        RECT 234.825 66.875 235.475 68.775 ;
        RECT 237.275 67.850 237.625 69.075 ;
        RECT 241.875 69.050 242.825 69.425 ;
        RECT 246.475 69.075 247.425 69.425 ;
        RECT 241.875 67.850 242.225 69.050 ;
        RECT 246.475 67.850 246.825 69.075 ;
        RECT 248.625 66.875 249.275 68.775 ;
        RECT 251.075 67.850 251.400 69.725 ;
        RECT 252.050 67.850 252.375 69.725 ;
        RECT 253.000 67.850 253.325 69.725 ;
        RECT 260.675 65.950 263.775 67.300 ;
        RECT 131.375 21.375 133.400 23.400 ;
        RECT 112.050 16.100 114.075 18.125 ;
        RECT 92.725 10.750 94.750 12.775 ;
        RECT 73.400 5.650 75.425 7.575 ;
      LAYER met3 ;
        RECT 126.450 215.100 127.600 217.150 ;
        RECT 138.275 213.850 139.100 214.450 ;
        RECT 135.525 210.575 136.350 211.175 ;
        RECT 132.775 207.300 133.600 207.900 ;
        RECT 130.000 204.050 130.825 204.650 ;
        RECT 111.925 200.575 113.050 201.100 ;
        RECT 180.125 200.575 181.250 201.100 ;
        RECT 68.000 195.850 73.160 199.250 ;
        RECT 76.490 195.850 81.650 199.250 ;
        RECT 84.980 195.850 90.140 199.250 ;
        RECT 93.470 195.850 98.630 199.250 ;
        RECT 101.960 195.850 107.120 199.250 ;
        RECT 110.000 195.850 115.160 199.250 ;
        RECT 118.490 195.850 123.650 199.250 ;
        RECT 126.980 195.850 132.140 199.250 ;
        RECT 135.470 195.850 140.630 199.250 ;
        RECT 143.960 195.850 149.120 199.250 ;
        RECT 152.000 195.850 157.160 199.250 ;
        RECT 160.490 195.850 165.650 199.250 ;
        RECT 168.980 195.850 174.140 199.250 ;
        RECT 177.010 195.850 182.170 199.250 ;
        RECT 185.500 195.850 190.660 199.250 ;
        RECT 193.990 195.850 199.150 199.250 ;
        RECT 202.000 195.850 207.160 199.250 ;
        RECT 210.000 195.850 215.160 199.250 ;
        RECT 68.000 190.850 73.160 194.250 ;
        RECT 76.490 190.850 81.650 194.250 ;
        RECT 84.980 190.850 90.140 194.250 ;
        RECT 93.470 190.850 98.630 194.250 ;
        RECT 101.960 190.850 107.120 194.250 ;
        RECT 110.000 190.850 115.160 194.250 ;
        RECT 118.490 190.850 123.650 194.250 ;
        RECT 126.980 190.850 132.140 194.250 ;
        RECT 135.470 190.850 140.630 194.250 ;
        RECT 143.960 190.850 149.120 194.250 ;
        RECT 152.000 190.850 157.160 194.250 ;
        RECT 160.490 190.850 165.650 194.250 ;
        RECT 168.980 190.850 174.140 194.250 ;
        RECT 177.010 190.850 182.170 194.250 ;
        RECT 185.500 190.850 190.660 194.250 ;
        RECT 193.990 190.850 199.150 194.250 ;
        RECT 202.000 190.850 207.160 194.250 ;
        RECT 210.000 190.850 215.160 194.250 ;
        RECT 68.000 185.850 73.160 189.250 ;
        RECT 76.490 185.850 81.650 189.250 ;
        RECT 84.980 185.850 90.140 189.250 ;
        RECT 93.470 185.850 98.630 189.250 ;
        RECT 101.960 185.850 107.120 189.250 ;
        RECT 110.000 185.850 115.160 189.250 ;
        RECT 118.490 185.850 123.650 189.250 ;
        RECT 126.980 185.850 132.140 189.250 ;
        RECT 135.470 185.850 140.630 189.250 ;
        RECT 143.960 185.850 149.120 189.250 ;
        RECT 152.000 185.850 157.160 189.250 ;
        RECT 160.490 185.850 165.650 189.250 ;
        RECT 168.980 185.850 174.140 189.250 ;
        RECT 177.010 185.850 182.170 189.250 ;
        RECT 185.500 185.850 190.660 189.250 ;
        RECT 193.990 185.850 199.150 189.250 ;
        RECT 202.000 185.850 207.160 189.250 ;
        RECT 210.000 185.850 215.160 189.250 ;
        RECT 68.000 180.850 73.160 184.250 ;
        RECT 76.490 180.850 81.650 184.250 ;
        RECT 84.980 180.850 90.140 184.250 ;
        RECT 93.470 180.850 98.630 184.250 ;
        RECT 101.960 180.850 107.120 184.250 ;
        RECT 110.000 180.850 115.160 184.250 ;
        RECT 118.490 180.850 123.650 184.250 ;
        RECT 126.980 180.850 132.140 184.250 ;
        RECT 135.470 180.850 140.630 184.250 ;
        RECT 143.960 180.850 149.120 184.250 ;
        RECT 152.000 180.850 157.160 184.250 ;
        RECT 160.490 180.850 165.650 184.250 ;
        RECT 168.980 180.850 174.140 184.250 ;
        RECT 177.010 180.850 182.170 184.250 ;
        RECT 185.500 180.850 190.660 184.250 ;
        RECT 193.990 180.850 199.150 184.250 ;
        RECT 202.000 180.850 207.160 184.250 ;
        RECT 210.000 180.850 215.160 184.250 ;
        RECT 68.000 175.850 73.160 179.250 ;
        RECT 76.490 175.850 81.650 179.250 ;
        RECT 84.980 175.850 90.140 179.250 ;
        RECT 93.470 175.850 98.630 179.250 ;
        RECT 101.960 175.850 107.120 179.250 ;
        RECT 110.000 175.850 115.160 179.250 ;
        RECT 118.490 175.850 123.650 179.250 ;
        RECT 126.980 175.850 132.140 179.250 ;
        RECT 135.470 175.850 140.630 179.250 ;
        RECT 143.960 175.850 149.120 179.250 ;
        RECT 152.000 175.850 157.160 179.250 ;
        RECT 160.490 175.850 165.650 179.250 ;
        RECT 168.980 175.850 174.140 179.250 ;
        RECT 177.010 175.850 182.170 179.250 ;
        RECT 185.500 175.850 190.660 179.250 ;
        RECT 193.990 175.850 199.150 179.250 ;
        RECT 202.000 175.850 207.160 179.250 ;
        RECT 210.000 175.850 215.160 179.250 ;
        RECT 68.000 170.850 73.160 174.250 ;
        RECT 76.490 170.850 81.650 174.250 ;
        RECT 84.980 170.850 90.140 174.250 ;
        RECT 93.470 170.850 98.630 174.250 ;
        RECT 101.960 170.850 107.120 174.250 ;
        RECT 110.000 170.850 115.160 174.250 ;
        RECT 118.490 170.850 123.650 174.250 ;
        RECT 126.980 170.850 132.140 174.250 ;
        RECT 135.470 170.850 140.630 174.250 ;
        RECT 143.960 170.850 149.120 174.250 ;
        RECT 152.000 170.850 157.160 174.250 ;
        RECT 160.490 170.850 165.650 174.250 ;
        RECT 168.980 170.850 174.140 174.250 ;
        RECT 177.010 170.850 182.170 174.250 ;
        RECT 185.500 170.850 190.660 174.250 ;
        RECT 193.990 170.850 199.150 174.250 ;
        RECT 68.000 165.850 73.160 169.250 ;
        RECT 76.490 165.850 81.650 169.250 ;
        RECT 84.980 165.850 90.140 169.250 ;
        RECT 93.470 165.850 98.630 169.250 ;
        RECT 101.960 165.850 107.120 169.250 ;
        RECT 110.000 165.850 115.160 169.250 ;
        RECT 118.490 165.850 123.650 169.250 ;
        RECT 126.980 165.850 132.140 169.250 ;
        RECT 135.470 165.850 140.630 169.250 ;
        RECT 143.960 165.850 149.120 169.250 ;
        RECT 152.000 165.850 157.160 169.250 ;
        RECT 160.490 165.850 165.650 169.250 ;
        RECT 168.980 165.850 174.140 169.250 ;
        RECT 177.010 165.850 182.170 169.250 ;
        RECT 185.500 165.850 190.660 169.250 ;
        RECT 193.990 165.850 199.150 169.250 ;
        RECT 65.000 129.375 71.000 149.900 ;
        RECT 1.000 123.450 71.000 129.375 ;
        RECT 4.000 104.275 59.700 110.200 ;
        RECT 65.000 94.675 71.000 123.450 ;
        RECT 72.650 82.500 73.525 137.250 ;
        RECT 75.275 67.675 81.175 158.225 ;
        RECT 203.125 154.850 204.250 173.325 ;
        RECT 206.200 163.200 259.050 164.275 ;
        RECT 179.225 153.725 204.250 154.850 ;
        RECT 212.800 161.250 259.050 163.200 ;
        RECT 179.225 153.150 180.350 153.725 ;
        RECT 122.000 151.425 180.350 153.150 ;
        RECT 122.000 150.720 124.050 151.425 ;
        RECT 212.800 150.720 215.825 161.250 ;
        RECT 240.925 158.275 246.250 159.000 ;
        RECT 84.605 148.670 124.055 150.720 ;
        RECT 84.605 135.845 86.655 148.670 ;
        RECT 98.030 141.820 112.680 143.370 ;
        RECT 90.725 127.200 91.850 133.775 ;
        RECT 97.930 130.670 99.980 137.395 ;
        RECT 122.005 135.845 124.055 148.670 ;
        RECT 135.330 148.670 215.830 150.720 ;
        RECT 135.330 141.820 136.880 148.670 ;
        RECT 161.980 141.820 163.530 148.670 ;
        RECT 128.605 138.270 190.055 139.820 ;
        RECT 128.605 134.645 130.155 138.270 ;
        RECT 122.105 133.095 130.155 134.645 ;
        RECT 135.330 130.670 137.380 137.395 ;
        RECT 148.655 135.845 150.705 138.270 ;
        RECT 161.980 135.845 164.030 138.270 ;
        RECT 97.930 128.620 137.380 130.670 ;
        RECT 148.655 130.670 150.205 134.645 ;
        RECT 173.705 130.670 175.755 137.620 ;
        RECT 176.380 135.320 178.430 137.395 ;
        RECT 189.705 135.320 191.755 137.395 ;
        RECT 199.380 135.845 201.430 148.670 ;
        RECT 212.805 141.820 227.455 143.370 ;
        RECT 206.005 135.845 213.155 137.395 ;
        RECT 206.005 135.320 207.555 135.845 ;
        RECT 176.380 133.770 207.555 135.320 ;
        RECT 213.780 130.675 215.830 137.395 ;
        RECT 212.800 130.670 215.830 130.675 ;
        RECT 148.655 128.620 215.830 130.670 ;
        RECT 135.325 127.950 137.375 128.620 ;
        RECT 90.725 126.075 113.050 127.200 ;
        RECT 135.325 126.225 211.350 127.950 ;
        RECT 88.700 118.725 93.860 122.125 ;
        RECT 97.190 118.725 102.350 122.125 ;
        RECT 105.680 118.725 110.840 122.125 ;
        RECT 114.170 118.725 119.330 122.125 ;
        RECT 122.660 118.725 127.820 122.125 ;
        RECT 131.150 118.725 136.310 122.125 ;
        RECT 139.640 118.725 144.800 122.125 ;
        RECT 148.130 118.725 153.290 122.125 ;
        RECT 156.620 118.725 161.780 122.125 ;
        RECT 165.110 118.725 170.270 122.125 ;
        RECT 173.600 118.725 178.760 122.125 ;
        RECT 182.090 118.725 187.250 122.125 ;
        RECT 190.580 118.725 195.740 122.125 ;
        RECT 199.070 118.725 204.230 122.125 ;
        RECT 206.450 122.025 207.800 124.150 ;
        RECT 212.800 118.050 215.825 128.620 ;
        RECT 234.375 120.300 235.925 152.500 ;
        RECT 238.975 124.750 240.525 157.900 ;
        RECT 240.925 153.975 241.650 158.275 ;
        RECT 240.925 153.375 241.975 153.975 ;
        RECT 240.925 145.875 241.650 153.375 ;
        RECT 242.450 149.750 243.175 153.975 ;
        RECT 240.925 145.150 243.050 145.875 ;
        RECT 243.575 145.600 245.125 157.900 ;
        RECT 245.525 153.975 246.250 158.275 ;
        RECT 245.525 153.375 246.575 153.975 ;
        RECT 242.450 144.675 243.050 145.150 ;
        RECT 246.100 144.675 246.825 150.400 ;
        RECT 240.925 144.075 241.975 144.675 ;
        RECT 242.450 144.075 243.175 144.675 ;
        RECT 245.775 144.075 246.825 144.675 ;
        RECT 240.925 143.600 241.650 144.075 ;
        RECT 246.100 143.600 246.825 144.075 ;
        RECT 240.925 142.875 246.825 143.600 ;
        RECT 240.925 137.425 246.250 138.150 ;
        RECT 240.925 133.125 241.650 137.425 ;
        RECT 240.925 132.525 241.975 133.125 ;
        RECT 240.925 125.025 241.650 132.525 ;
        RECT 242.450 128.900 243.175 133.125 ;
        RECT 240.925 124.300 243.050 125.025 ;
        RECT 243.575 124.750 245.125 137.050 ;
        RECT 245.525 133.125 246.250 137.425 ;
        RECT 245.525 132.525 246.575 133.125 ;
        RECT 242.450 123.825 243.050 124.300 ;
        RECT 246.100 123.825 246.825 129.550 ;
        RECT 240.925 123.225 241.975 123.825 ;
        RECT 242.450 123.225 243.175 123.825 ;
        RECT 245.775 123.225 246.825 123.825 ;
        RECT 240.925 122.750 241.650 123.225 ;
        RECT 246.100 122.750 246.825 123.225 ;
        RECT 240.925 122.025 246.825 122.750 ;
        RECT 248.175 120.300 249.725 152.500 ;
        RECT 254.950 145.750 259.050 161.250 ;
        RECT 258.350 135.950 261.450 141.650 ;
        RECT 263.300 137.650 266.400 159.850 ;
        RECT 258.350 132.850 263.775 135.950 ;
        RECT 254.950 118.050 259.050 131.275 ;
        RECT 260.675 119.450 263.775 132.850 ;
        RECT 88.700 113.725 93.860 117.125 ;
        RECT 97.190 113.725 102.350 117.125 ;
        RECT 105.680 113.725 110.840 117.125 ;
        RECT 114.170 113.725 119.330 117.125 ;
        RECT 122.660 113.725 127.820 117.125 ;
        RECT 131.150 113.725 136.310 117.125 ;
        RECT 139.640 113.725 144.800 117.125 ;
        RECT 148.130 113.725 153.290 117.125 ;
        RECT 156.620 113.725 161.780 117.125 ;
        RECT 165.110 113.725 170.270 117.125 ;
        RECT 173.600 113.725 178.760 117.125 ;
        RECT 182.090 113.725 187.250 117.125 ;
        RECT 190.580 113.725 195.740 117.125 ;
        RECT 199.070 113.725 204.230 117.125 ;
        RECT 212.800 115.000 259.050 118.050 ;
        RECT 88.700 108.725 93.860 112.125 ;
        RECT 97.190 108.725 102.350 112.125 ;
        RECT 105.680 108.725 110.840 112.125 ;
        RECT 114.170 108.725 119.330 112.125 ;
        RECT 122.660 108.725 127.820 112.125 ;
        RECT 131.150 108.725 136.310 112.125 ;
        RECT 139.640 108.725 144.800 112.125 ;
        RECT 148.130 108.725 153.290 112.125 ;
        RECT 156.620 108.725 161.780 112.125 ;
        RECT 165.110 108.725 170.270 112.125 ;
        RECT 173.600 108.725 178.760 112.125 ;
        RECT 182.090 108.725 187.250 112.125 ;
        RECT 190.580 108.725 195.740 112.125 ;
        RECT 199.070 108.725 204.230 112.125 ;
        RECT 212.800 107.750 259.050 110.775 ;
        RECT 88.700 103.725 93.860 107.125 ;
        RECT 97.190 103.725 102.350 107.125 ;
        RECT 105.680 103.725 110.840 107.125 ;
        RECT 114.170 103.725 119.330 107.125 ;
        RECT 122.660 103.725 127.820 107.125 ;
        RECT 131.150 103.725 136.310 107.125 ;
        RECT 139.640 103.725 144.800 107.125 ;
        RECT 148.130 103.725 153.290 107.125 ;
        RECT 156.620 103.725 161.780 107.125 ;
        RECT 165.110 103.725 170.270 107.125 ;
        RECT 173.600 103.725 178.760 107.125 ;
        RECT 182.090 103.725 187.250 107.125 ;
        RECT 190.580 103.725 195.740 107.125 ;
        RECT 199.070 103.725 204.230 107.125 ;
        RECT 206.450 101.750 207.800 103.825 ;
        RECT 82.400 98.775 113.050 99.825 ;
        RECT 82.400 91.900 83.525 98.775 ;
        RECT 122.000 97.925 211.350 99.650 ;
        RECT 122.000 97.220 124.050 97.925 ;
        RECT 212.800 97.220 215.825 107.750 ;
        RECT 240.925 104.775 246.250 105.500 ;
        RECT 84.605 95.170 124.055 97.220 ;
        RECT 84.605 82.345 86.655 95.170 ;
        RECT 98.030 88.320 112.680 89.870 ;
        RECT 97.930 77.170 99.980 83.895 ;
        RECT 122.005 82.345 124.055 95.170 ;
        RECT 135.330 95.170 215.830 97.220 ;
        RECT 135.330 88.320 136.880 95.170 ;
        RECT 161.980 88.320 163.530 95.170 ;
        RECT 128.605 84.770 190.055 86.320 ;
        RECT 128.605 81.145 130.155 84.770 ;
        RECT 122.105 79.595 130.155 81.145 ;
        RECT 135.330 77.170 137.380 83.895 ;
        RECT 148.655 82.345 150.705 84.770 ;
        RECT 161.980 82.345 164.030 84.770 ;
        RECT 97.930 75.120 137.380 77.170 ;
        RECT 148.655 77.170 150.205 81.145 ;
        RECT 173.705 77.170 175.755 84.120 ;
        RECT 176.380 81.820 178.430 83.895 ;
        RECT 189.705 81.820 191.755 83.895 ;
        RECT 199.380 82.345 201.430 95.170 ;
        RECT 212.805 88.320 227.455 89.870 ;
        RECT 206.005 82.345 213.155 83.895 ;
        RECT 206.005 81.820 207.555 82.345 ;
        RECT 176.380 80.270 207.555 81.820 ;
        RECT 213.780 77.175 215.830 83.895 ;
        RECT 212.800 77.170 215.830 77.175 ;
        RECT 148.655 75.120 215.830 77.170 ;
        RECT 135.325 74.450 137.375 75.120 ;
        RECT 135.325 72.725 180.350 74.450 ;
        RECT 179.225 72.150 180.350 72.725 ;
        RECT 179.225 71.025 204.250 72.150 ;
        RECT 68.000 56.850 73.160 60.250 ;
        RECT 76.490 56.850 81.650 60.250 ;
        RECT 84.980 56.850 90.140 60.250 ;
        RECT 93.470 56.850 98.630 60.250 ;
        RECT 101.960 56.850 107.120 60.250 ;
        RECT 110.000 56.850 115.160 60.250 ;
        RECT 118.490 56.850 123.650 60.250 ;
        RECT 126.980 56.850 132.140 60.250 ;
        RECT 135.470 56.850 140.630 60.250 ;
        RECT 143.960 56.850 149.120 60.250 ;
        RECT 152.000 56.850 157.160 60.250 ;
        RECT 160.490 56.850 165.650 60.250 ;
        RECT 168.980 56.850 174.140 60.250 ;
        RECT 177.010 56.850 182.170 60.250 ;
        RECT 185.500 56.850 190.660 60.250 ;
        RECT 193.990 56.850 199.150 60.250 ;
        RECT 68.000 51.850 73.160 55.250 ;
        RECT 76.490 51.850 81.650 55.250 ;
        RECT 84.980 51.850 90.140 55.250 ;
        RECT 93.470 51.850 98.630 55.250 ;
        RECT 101.960 51.850 107.120 55.250 ;
        RECT 110.000 51.850 115.160 55.250 ;
        RECT 118.490 51.850 123.650 55.250 ;
        RECT 126.980 51.850 132.140 55.250 ;
        RECT 135.470 51.850 140.630 55.250 ;
        RECT 143.960 51.850 149.120 55.250 ;
        RECT 152.000 51.850 157.160 55.250 ;
        RECT 160.490 51.850 165.650 55.250 ;
        RECT 168.980 51.850 174.140 55.250 ;
        RECT 177.010 51.850 182.170 55.250 ;
        RECT 185.500 51.850 190.660 55.250 ;
        RECT 193.990 51.850 199.150 55.250 ;
        RECT 203.125 52.550 204.250 71.025 ;
        RECT 212.800 64.550 215.825 75.120 ;
        RECT 234.375 66.800 235.925 99.000 ;
        RECT 238.975 71.250 240.525 104.400 ;
        RECT 240.925 100.475 241.650 104.775 ;
        RECT 240.925 99.875 241.975 100.475 ;
        RECT 240.925 92.375 241.650 99.875 ;
        RECT 242.450 96.250 243.175 100.475 ;
        RECT 240.925 91.650 243.050 92.375 ;
        RECT 243.575 92.100 245.125 104.400 ;
        RECT 245.525 100.475 246.250 104.775 ;
        RECT 245.525 99.875 246.575 100.475 ;
        RECT 242.450 91.175 243.050 91.650 ;
        RECT 246.100 91.175 246.825 96.900 ;
        RECT 240.925 90.575 241.975 91.175 ;
        RECT 242.450 90.575 243.175 91.175 ;
        RECT 245.775 90.575 246.825 91.175 ;
        RECT 240.925 90.100 241.650 90.575 ;
        RECT 246.100 90.100 246.825 90.575 ;
        RECT 240.925 89.375 246.825 90.100 ;
        RECT 240.925 83.925 246.250 84.650 ;
        RECT 240.925 79.625 241.650 83.925 ;
        RECT 240.925 79.025 241.975 79.625 ;
        RECT 240.925 71.525 241.650 79.025 ;
        RECT 242.450 75.400 243.175 79.625 ;
        RECT 240.925 70.800 243.050 71.525 ;
        RECT 243.575 71.250 245.125 83.550 ;
        RECT 245.525 79.625 246.250 83.925 ;
        RECT 245.525 79.025 246.575 79.625 ;
        RECT 242.450 70.325 243.050 70.800 ;
        RECT 246.100 70.325 246.825 76.050 ;
        RECT 240.925 69.725 241.975 70.325 ;
        RECT 242.450 69.725 243.175 70.325 ;
        RECT 245.775 69.725 246.825 70.325 ;
        RECT 240.925 69.250 241.650 69.725 ;
        RECT 246.100 69.250 246.825 69.725 ;
        RECT 240.925 68.525 246.825 69.250 ;
        RECT 248.175 66.800 249.725 99.000 ;
        RECT 254.950 92.250 259.050 107.750 ;
        RECT 265.075 106.350 266.400 137.650 ;
        RECT 268.350 124.900 275.150 152.125 ;
        RECT 258.350 82.450 261.450 88.150 ;
        RECT 263.300 84.150 266.400 106.350 ;
        RECT 270.600 98.625 275.150 124.900 ;
        RECT 258.350 79.350 263.775 82.450 ;
        RECT 254.950 64.550 259.050 77.775 ;
        RECT 260.675 65.950 263.775 79.350 ;
        RECT 268.350 71.400 275.150 98.625 ;
        RECT 212.800 62.575 259.050 64.550 ;
        RECT 206.225 61.500 259.050 62.575 ;
        RECT 68.000 46.850 73.160 50.250 ;
        RECT 76.490 46.850 81.650 50.250 ;
        RECT 84.980 46.850 90.140 50.250 ;
        RECT 93.470 46.850 98.630 50.250 ;
        RECT 101.960 46.850 107.120 50.250 ;
        RECT 110.000 46.850 115.160 50.250 ;
        RECT 118.490 46.850 123.650 50.250 ;
        RECT 126.980 46.850 132.140 50.250 ;
        RECT 135.470 46.850 140.630 50.250 ;
        RECT 143.960 46.850 149.120 50.250 ;
        RECT 152.000 46.850 157.160 50.250 ;
        RECT 160.490 46.850 165.650 50.250 ;
        RECT 168.980 46.850 174.140 50.250 ;
        RECT 177.010 46.850 182.170 50.250 ;
        RECT 185.500 46.850 190.660 50.250 ;
        RECT 193.990 46.850 199.150 50.250 ;
        RECT 202.000 46.850 207.160 50.250 ;
        RECT 210.000 46.850 215.160 50.250 ;
        RECT 68.000 41.850 73.160 45.250 ;
        RECT 76.490 41.850 81.650 45.250 ;
        RECT 84.980 41.850 90.140 45.250 ;
        RECT 93.470 41.850 98.630 45.250 ;
        RECT 101.960 41.850 107.120 45.250 ;
        RECT 110.000 41.850 115.160 45.250 ;
        RECT 118.490 41.850 123.650 45.250 ;
        RECT 126.980 41.850 132.140 45.250 ;
        RECT 135.470 41.850 140.630 45.250 ;
        RECT 143.960 41.850 149.120 45.250 ;
        RECT 152.000 41.850 157.160 45.250 ;
        RECT 160.490 41.850 165.650 45.250 ;
        RECT 168.980 41.850 174.140 45.250 ;
        RECT 177.010 41.850 182.170 45.250 ;
        RECT 185.500 41.850 190.660 45.250 ;
        RECT 193.990 41.850 199.150 45.250 ;
        RECT 202.000 41.850 207.160 45.250 ;
        RECT 210.000 41.850 215.160 45.250 ;
        RECT 68.000 36.850 73.160 40.250 ;
        RECT 76.490 36.850 81.650 40.250 ;
        RECT 84.980 36.850 90.140 40.250 ;
        RECT 93.470 36.850 98.630 40.250 ;
        RECT 101.960 36.850 107.120 40.250 ;
        RECT 110.000 36.850 115.160 40.250 ;
        RECT 118.490 36.850 123.650 40.250 ;
        RECT 126.980 36.850 132.140 40.250 ;
        RECT 135.470 36.850 140.630 40.250 ;
        RECT 143.960 36.850 149.120 40.250 ;
        RECT 152.000 36.850 157.160 40.250 ;
        RECT 160.490 36.850 165.650 40.250 ;
        RECT 168.980 36.850 174.140 40.250 ;
        RECT 177.010 36.850 182.170 40.250 ;
        RECT 185.500 36.850 190.660 40.250 ;
        RECT 193.990 36.850 199.150 40.250 ;
        RECT 202.000 36.850 207.160 40.250 ;
        RECT 210.000 36.850 215.160 40.250 ;
        RECT 68.000 31.850 73.160 35.250 ;
        RECT 76.490 31.850 81.650 35.250 ;
        RECT 84.980 31.850 90.140 35.250 ;
        RECT 93.470 31.850 98.630 35.250 ;
        RECT 101.960 31.850 107.120 35.250 ;
        RECT 110.000 31.850 115.160 35.250 ;
        RECT 118.490 31.850 123.650 35.250 ;
        RECT 126.980 31.850 132.140 35.250 ;
        RECT 135.470 31.850 140.630 35.250 ;
        RECT 143.960 31.850 149.120 35.250 ;
        RECT 152.000 31.850 157.160 35.250 ;
        RECT 160.490 31.850 165.650 35.250 ;
        RECT 168.980 31.850 174.140 35.250 ;
        RECT 177.010 31.850 182.170 35.250 ;
        RECT 185.500 31.850 190.660 35.250 ;
        RECT 193.990 31.850 199.150 35.250 ;
        RECT 202.000 31.850 207.160 35.250 ;
        RECT 210.000 31.850 215.160 35.250 ;
        RECT 68.000 26.850 73.160 30.250 ;
        RECT 76.490 26.850 81.650 30.250 ;
        RECT 84.980 26.850 90.140 30.250 ;
        RECT 93.470 26.850 98.630 30.250 ;
        RECT 101.960 26.850 107.120 30.250 ;
        RECT 110.000 26.850 115.160 30.250 ;
        RECT 118.490 26.850 123.650 30.250 ;
        RECT 126.980 26.850 132.140 30.250 ;
        RECT 135.470 26.850 140.630 30.250 ;
        RECT 143.960 26.850 149.120 30.250 ;
        RECT 152.000 26.850 157.160 30.250 ;
        RECT 160.490 26.850 165.650 30.250 ;
        RECT 168.980 26.850 174.140 30.250 ;
        RECT 177.010 26.850 182.170 30.250 ;
        RECT 185.500 26.850 190.660 30.250 ;
        RECT 193.990 26.850 199.150 30.250 ;
        RECT 202.000 26.850 207.160 30.250 ;
        RECT 210.000 26.850 215.160 30.250 ;
        RECT 111.925 25.000 113.050 25.525 ;
        RECT 180.125 25.000 181.250 25.525 ;
        RECT 131.375 21.375 133.400 23.400 ;
        RECT 112.050 16.100 114.075 18.125 ;
        RECT 92.725 10.750 94.750 12.775 ;
        RECT 272.100 8.700 275.150 71.400 ;
        RECT 73.400 5.650 75.425 7.575 ;
        RECT 151.800 5.650 275.150 8.700 ;
      LAYER met4 ;
        RECT 127.250 224.760 127.270 225.300 ;
        RECT 127.570 224.760 127.600 225.300 ;
        RECT 127.250 217.150 127.600 224.760 ;
        RECT 126.450 215.100 127.600 217.150 ;
        RECT 130.000 224.760 130.030 225.300 ;
        RECT 130.330 224.760 130.350 225.300 ;
        RECT 130.000 204.650 130.350 224.760 ;
        RECT 132.775 224.760 132.790 225.300 ;
        RECT 133.090 224.760 133.125 225.300 ;
        RECT 132.775 207.900 133.125 224.760 ;
        RECT 135.525 224.760 135.550 225.300 ;
        RECT 135.850 224.760 135.875 225.300 ;
        RECT 135.525 211.175 135.875 224.760 ;
        RECT 138.275 224.760 138.310 225.300 ;
        RECT 138.610 224.760 138.625 225.300 ;
        RECT 138.275 214.450 138.625 224.760 ;
        RECT 138.275 213.850 139.100 214.450 ;
        RECT 135.525 210.575 136.350 211.175 ;
        RECT 132.775 207.300 133.600 207.900 ;
        RECT 130.000 204.050 130.825 204.650 ;
        RECT 69.435 200.575 144.485 201.100 ;
        RECT 69.435 200.050 69.960 200.575 ;
        RECT 77.935 200.050 78.460 200.575 ;
        RECT 86.410 200.050 86.935 200.575 ;
        RECT 94.910 200.050 95.435 200.575 ;
        RECT 103.385 200.050 103.910 200.575 ;
        RECT 110.010 200.050 110.535 200.575 ;
        RECT 118.485 200.050 119.010 200.575 ;
        RECT 126.985 200.050 127.510 200.575 ;
        RECT 135.460 200.050 135.985 200.575 ;
        RECT 143.960 200.050 144.485 200.575 ;
        RECT 153.450 200.575 194.500 201.100 ;
        RECT 203.400 200.575 203.975 201.100 ;
        RECT 211.400 200.575 211.975 201.100 ;
        RECT 153.450 200.050 153.975 200.575 ;
        RECT 161.950 200.050 162.475 200.575 ;
        RECT 170.425 200.050 170.950 200.575 ;
        RECT 177.000 200.050 177.525 200.575 ;
        RECT 185.475 200.050 186.000 200.575 ;
        RECT 193.975 200.050 194.500 200.575 ;
        RECT 203.425 200.050 203.950 200.575 ;
        RECT 211.425 200.050 211.950 200.575 ;
        RECT 69.440 198.855 69.960 200.050 ;
        RECT 68.395 196.245 71.005 198.855 ;
        RECT 69.440 193.855 69.960 196.245 ;
        RECT 68.395 191.245 71.005 193.855 ;
        RECT 69.440 188.855 69.960 191.245 ;
        RECT 68.395 186.245 71.005 188.855 ;
        RECT 69.440 183.855 69.960 186.245 ;
        RECT 68.395 181.245 71.005 183.855 ;
        RECT 69.440 178.855 69.960 181.245 ;
        RECT 68.395 176.245 71.005 178.855 ;
        RECT 69.440 173.855 69.960 176.245 ;
        RECT 68.395 171.245 71.005 173.855 ;
        RECT 69.440 168.855 69.960 171.245 ;
        RECT 68.395 166.245 71.005 168.855 ;
        RECT 69.440 165.050 69.960 166.245 ;
        RECT 72.640 165.050 73.160 200.050 ;
        RECT 77.930 198.855 78.450 200.050 ;
        RECT 76.885 196.245 79.495 198.855 ;
        RECT 77.930 193.855 78.450 196.245 ;
        RECT 76.885 191.245 79.495 193.855 ;
        RECT 77.930 188.855 78.450 191.245 ;
        RECT 76.885 186.245 79.495 188.855 ;
        RECT 77.930 183.855 78.450 186.245 ;
        RECT 76.885 181.245 79.495 183.855 ;
        RECT 77.930 178.855 78.450 181.245 ;
        RECT 76.885 176.245 79.495 178.855 ;
        RECT 77.930 173.855 78.450 176.245 ;
        RECT 76.885 171.245 79.495 173.855 ;
        RECT 77.930 168.855 78.450 171.245 ;
        RECT 76.885 166.245 79.495 168.855 ;
        RECT 77.930 165.050 78.450 166.245 ;
        RECT 81.130 165.050 81.650 200.050 ;
        RECT 86.420 198.855 86.940 200.050 ;
        RECT 85.375 196.245 87.985 198.855 ;
        RECT 86.420 193.855 86.940 196.245 ;
        RECT 85.375 191.245 87.985 193.855 ;
        RECT 86.420 188.855 86.940 191.245 ;
        RECT 85.375 186.245 87.985 188.855 ;
        RECT 86.420 183.855 86.940 186.245 ;
        RECT 85.375 181.245 87.985 183.855 ;
        RECT 86.420 178.855 86.940 181.245 ;
        RECT 85.375 176.245 87.985 178.855 ;
        RECT 86.420 173.855 86.940 176.245 ;
        RECT 85.375 171.245 87.985 173.855 ;
        RECT 86.420 168.855 86.940 171.245 ;
        RECT 85.375 166.245 87.985 168.855 ;
        RECT 86.420 165.050 86.940 166.245 ;
        RECT 89.620 165.050 90.140 200.050 ;
        RECT 94.910 198.855 95.430 200.050 ;
        RECT 93.865 196.245 96.475 198.855 ;
        RECT 94.910 193.855 95.430 196.245 ;
        RECT 93.865 191.245 96.475 193.855 ;
        RECT 94.910 188.855 95.430 191.245 ;
        RECT 93.865 186.245 96.475 188.855 ;
        RECT 94.910 183.855 95.430 186.245 ;
        RECT 93.865 181.245 96.475 183.855 ;
        RECT 94.910 178.855 95.430 181.245 ;
        RECT 93.865 176.245 96.475 178.855 ;
        RECT 94.910 173.855 95.430 176.245 ;
        RECT 93.865 171.245 96.475 173.855 ;
        RECT 94.910 168.855 95.430 171.245 ;
        RECT 93.865 166.245 96.475 168.855 ;
        RECT 94.910 165.050 95.430 166.245 ;
        RECT 98.110 165.050 98.630 200.050 ;
        RECT 103.400 198.855 103.920 200.050 ;
        RECT 102.355 196.245 104.965 198.855 ;
        RECT 103.400 193.855 103.920 196.245 ;
        RECT 102.355 191.245 104.965 193.855 ;
        RECT 103.400 188.855 103.920 191.245 ;
        RECT 102.355 186.245 104.965 188.855 ;
        RECT 103.400 183.855 103.920 186.245 ;
        RECT 102.355 181.245 104.965 183.855 ;
        RECT 103.400 178.855 103.920 181.245 ;
        RECT 102.355 176.245 104.965 178.855 ;
        RECT 103.400 173.855 103.920 176.245 ;
        RECT 102.355 171.245 104.965 173.855 ;
        RECT 103.400 168.855 103.920 171.245 ;
        RECT 102.355 166.245 104.965 168.855 ;
        RECT 103.400 165.050 103.920 166.245 ;
        RECT 106.600 165.050 107.120 200.050 ;
        RECT 110.000 165.050 110.520 200.050 ;
        RECT 113.200 198.855 113.720 200.050 ;
        RECT 112.155 196.245 114.765 198.855 ;
        RECT 113.200 193.855 113.720 196.245 ;
        RECT 112.155 191.245 114.765 193.855 ;
        RECT 113.200 188.855 113.720 191.245 ;
        RECT 112.155 186.245 114.765 188.855 ;
        RECT 113.200 183.855 113.720 186.245 ;
        RECT 112.155 181.245 114.765 183.855 ;
        RECT 113.200 178.855 113.720 181.245 ;
        RECT 112.155 176.245 114.765 178.855 ;
        RECT 113.200 173.855 113.720 176.245 ;
        RECT 112.155 171.245 114.765 173.855 ;
        RECT 113.200 168.855 113.720 171.245 ;
        RECT 112.155 166.245 114.765 168.855 ;
        RECT 113.200 165.050 113.720 166.245 ;
        RECT 118.490 165.050 119.010 200.050 ;
        RECT 121.690 198.855 122.210 200.050 ;
        RECT 120.645 196.245 123.255 198.855 ;
        RECT 121.690 193.855 122.210 196.245 ;
        RECT 120.645 191.245 123.255 193.855 ;
        RECT 121.690 188.855 122.210 191.245 ;
        RECT 120.645 186.245 123.255 188.855 ;
        RECT 121.690 183.855 122.210 186.245 ;
        RECT 120.645 181.245 123.255 183.855 ;
        RECT 121.690 178.855 122.210 181.245 ;
        RECT 120.645 176.245 123.255 178.855 ;
        RECT 121.690 173.855 122.210 176.245 ;
        RECT 120.645 171.245 123.255 173.855 ;
        RECT 121.690 168.855 122.210 171.245 ;
        RECT 120.645 166.245 123.255 168.855 ;
        RECT 121.690 165.050 122.210 166.245 ;
        RECT 126.980 165.050 127.500 200.050 ;
        RECT 130.180 198.855 130.700 200.050 ;
        RECT 129.135 196.245 131.745 198.855 ;
        RECT 130.180 193.855 130.700 196.245 ;
        RECT 129.135 191.245 131.745 193.855 ;
        RECT 130.180 188.855 130.700 191.245 ;
        RECT 129.135 186.245 131.745 188.855 ;
        RECT 130.180 183.855 130.700 186.245 ;
        RECT 129.135 181.245 131.745 183.855 ;
        RECT 130.180 178.855 130.700 181.245 ;
        RECT 129.135 176.245 131.745 178.855 ;
        RECT 130.180 173.855 130.700 176.245 ;
        RECT 129.135 171.245 131.745 173.855 ;
        RECT 130.180 168.855 130.700 171.245 ;
        RECT 129.135 166.245 131.745 168.855 ;
        RECT 130.180 165.050 130.700 166.245 ;
        RECT 135.470 165.050 135.990 200.050 ;
        RECT 138.670 198.855 139.190 200.050 ;
        RECT 137.625 196.245 140.235 198.855 ;
        RECT 138.670 193.855 139.190 196.245 ;
        RECT 137.625 191.245 140.235 193.855 ;
        RECT 138.670 188.855 139.190 191.245 ;
        RECT 137.625 186.245 140.235 188.855 ;
        RECT 138.670 183.855 139.190 186.245 ;
        RECT 137.625 181.245 140.235 183.855 ;
        RECT 138.670 178.855 139.190 181.245 ;
        RECT 137.625 176.245 140.235 178.855 ;
        RECT 138.670 173.855 139.190 176.245 ;
        RECT 137.625 171.245 140.235 173.855 ;
        RECT 138.670 168.855 139.190 171.245 ;
        RECT 137.625 166.245 140.235 168.855 ;
        RECT 138.670 165.050 139.190 166.245 ;
        RECT 143.960 165.050 144.480 200.050 ;
        RECT 147.160 198.855 147.680 200.050 ;
        RECT 153.440 198.855 153.960 200.050 ;
        RECT 146.115 196.245 148.725 198.855 ;
        RECT 152.395 196.245 155.005 198.855 ;
        RECT 147.160 193.855 147.680 196.245 ;
        RECT 153.440 193.855 153.960 196.245 ;
        RECT 146.115 191.245 148.725 193.855 ;
        RECT 152.395 191.245 155.005 193.855 ;
        RECT 147.160 188.855 147.680 191.245 ;
        RECT 153.440 188.855 153.960 191.245 ;
        RECT 146.115 186.245 148.725 188.855 ;
        RECT 152.395 186.245 155.005 188.855 ;
        RECT 147.160 183.855 147.680 186.245 ;
        RECT 153.440 183.855 153.960 186.245 ;
        RECT 146.115 181.245 148.725 183.855 ;
        RECT 152.395 181.245 155.005 183.855 ;
        RECT 147.160 178.855 147.680 181.245 ;
        RECT 153.440 178.855 153.960 181.245 ;
        RECT 146.115 176.245 148.725 178.855 ;
        RECT 152.395 176.245 155.005 178.855 ;
        RECT 147.160 173.855 147.680 176.245 ;
        RECT 153.440 173.855 153.960 176.245 ;
        RECT 146.115 171.245 148.725 173.855 ;
        RECT 152.395 171.245 155.005 173.855 ;
        RECT 147.160 168.855 147.680 171.245 ;
        RECT 153.440 168.855 153.960 171.245 ;
        RECT 146.115 166.245 148.725 168.855 ;
        RECT 152.395 166.245 155.005 168.855 ;
        RECT 147.160 165.050 147.680 166.245 ;
        RECT 153.440 165.050 153.960 166.245 ;
        RECT 156.640 165.050 157.160 200.050 ;
        RECT 161.930 198.855 162.450 200.050 ;
        RECT 160.885 196.245 163.495 198.855 ;
        RECT 161.930 193.855 162.450 196.245 ;
        RECT 160.885 191.245 163.495 193.855 ;
        RECT 161.930 188.855 162.450 191.245 ;
        RECT 160.885 186.245 163.495 188.855 ;
        RECT 161.930 183.855 162.450 186.245 ;
        RECT 160.885 181.245 163.495 183.855 ;
        RECT 161.930 178.855 162.450 181.245 ;
        RECT 160.885 176.245 163.495 178.855 ;
        RECT 161.930 173.855 162.450 176.245 ;
        RECT 160.885 171.245 163.495 173.855 ;
        RECT 161.930 168.855 162.450 171.245 ;
        RECT 160.885 166.245 163.495 168.855 ;
        RECT 161.930 165.050 162.450 166.245 ;
        RECT 165.130 165.050 165.650 200.050 ;
        RECT 170.420 198.855 170.940 200.050 ;
        RECT 169.375 196.245 171.985 198.855 ;
        RECT 170.420 193.855 170.940 196.245 ;
        RECT 169.375 191.245 171.985 193.855 ;
        RECT 170.420 188.855 170.940 191.245 ;
        RECT 169.375 186.245 171.985 188.855 ;
        RECT 170.420 183.855 170.940 186.245 ;
        RECT 169.375 181.245 171.985 183.855 ;
        RECT 170.420 178.855 170.940 181.245 ;
        RECT 169.375 176.245 171.985 178.855 ;
        RECT 170.420 173.855 170.940 176.245 ;
        RECT 169.375 171.245 171.985 173.855 ;
        RECT 170.420 168.855 170.940 171.245 ;
        RECT 169.375 166.245 171.985 168.855 ;
        RECT 170.420 165.050 170.940 166.245 ;
        RECT 173.620 165.050 174.140 200.050 ;
        RECT 177.010 165.050 177.530 200.050 ;
        RECT 180.210 198.855 180.730 200.050 ;
        RECT 179.165 196.245 181.775 198.855 ;
        RECT 180.210 193.855 180.730 196.245 ;
        RECT 179.165 191.245 181.775 193.855 ;
        RECT 180.210 188.855 180.730 191.245 ;
        RECT 179.165 186.245 181.775 188.855 ;
        RECT 180.210 183.855 180.730 186.245 ;
        RECT 179.165 181.245 181.775 183.855 ;
        RECT 180.210 178.855 180.730 181.245 ;
        RECT 179.165 176.245 181.775 178.855 ;
        RECT 180.210 173.855 180.730 176.245 ;
        RECT 179.165 171.245 181.775 173.855 ;
        RECT 180.210 168.855 180.730 171.245 ;
        RECT 179.165 166.245 181.775 168.855 ;
        RECT 180.210 165.050 180.730 166.245 ;
        RECT 185.500 165.050 186.020 200.050 ;
        RECT 188.700 198.855 189.220 200.050 ;
        RECT 187.655 196.245 190.265 198.855 ;
        RECT 188.700 193.855 189.220 196.245 ;
        RECT 187.655 191.245 190.265 193.855 ;
        RECT 188.700 188.855 189.220 191.245 ;
        RECT 187.655 186.245 190.265 188.855 ;
        RECT 188.700 183.855 189.220 186.245 ;
        RECT 187.655 181.245 190.265 183.855 ;
        RECT 188.700 178.855 189.220 181.245 ;
        RECT 187.655 176.245 190.265 178.855 ;
        RECT 188.700 173.855 189.220 176.245 ;
        RECT 187.655 171.245 190.265 173.855 ;
        RECT 188.700 168.855 189.220 171.245 ;
        RECT 187.655 166.245 190.265 168.855 ;
        RECT 188.700 165.050 189.220 166.245 ;
        RECT 193.990 165.050 194.510 200.050 ;
        RECT 197.190 198.855 197.710 200.050 ;
        RECT 203.440 198.855 203.960 200.050 ;
        RECT 196.145 196.245 198.755 198.855 ;
        RECT 202.395 196.245 205.005 198.855 ;
        RECT 197.190 193.855 197.710 196.245 ;
        RECT 203.440 193.855 203.960 196.245 ;
        RECT 196.145 191.245 198.755 193.855 ;
        RECT 202.395 191.245 205.005 193.855 ;
        RECT 197.190 188.855 197.710 191.245 ;
        RECT 203.440 188.855 203.960 191.245 ;
        RECT 196.145 186.245 198.755 188.855 ;
        RECT 202.395 186.245 205.005 188.855 ;
        RECT 197.190 183.855 197.710 186.245 ;
        RECT 203.440 183.855 203.960 186.245 ;
        RECT 196.145 181.245 198.755 183.855 ;
        RECT 202.395 181.245 205.005 183.855 ;
        RECT 197.190 178.855 197.710 181.245 ;
        RECT 203.440 178.855 203.960 181.245 ;
        RECT 196.145 176.245 198.755 178.855 ;
        RECT 202.395 176.245 205.005 178.855 ;
        RECT 197.190 173.855 197.710 176.245 ;
        RECT 203.440 175.075 203.960 176.245 ;
        RECT 203.425 175.050 203.960 175.075 ;
        RECT 206.640 175.050 207.160 200.050 ;
        RECT 211.440 198.855 211.960 200.050 ;
        RECT 210.395 196.245 213.005 198.855 ;
        RECT 211.440 193.855 211.960 196.245 ;
        RECT 210.395 191.245 213.005 193.855 ;
        RECT 211.440 188.855 211.960 191.245 ;
        RECT 210.395 186.245 213.005 188.855 ;
        RECT 211.440 183.855 211.960 186.245 ;
        RECT 210.395 181.245 213.005 183.855 ;
        RECT 211.440 178.855 211.960 181.245 ;
        RECT 210.395 176.245 213.005 178.855 ;
        RECT 211.440 175.050 211.960 176.245 ;
        RECT 214.640 175.050 215.160 200.050 ;
        RECT 196.145 171.245 198.755 173.855 ;
        RECT 203.425 173.325 203.950 175.050 ;
        RECT 206.625 174.525 207.150 175.050 ;
        RECT 210.000 174.675 211.950 175.050 ;
        RECT 206.600 174.025 207.175 174.525 ;
        RECT 203.125 172.600 204.250 173.325 ;
        RECT 197.190 168.855 197.710 171.245 ;
        RECT 196.145 166.245 198.755 168.855 ;
        RECT 197.190 165.050 197.710 166.245 ;
        RECT 72.635 164.525 73.160 165.050 ;
        RECT 81.135 164.525 81.660 165.050 ;
        RECT 89.610 164.525 90.135 165.050 ;
        RECT 98.110 164.525 98.635 165.050 ;
        RECT 106.585 164.525 107.110 165.050 ;
        RECT 113.210 164.525 113.735 165.050 ;
        RECT 121.685 164.525 122.210 165.050 ;
        RECT 130.185 164.525 130.710 165.050 ;
        RECT 138.660 164.525 139.185 165.050 ;
        RECT 147.160 164.525 147.685 165.050 ;
        RECT 72.635 164.000 147.685 164.525 ;
        RECT 156.650 164.525 157.175 165.050 ;
        RECT 165.150 164.525 165.675 165.050 ;
        RECT 173.625 164.525 174.150 165.050 ;
        RECT 180.200 164.525 180.725 165.050 ;
        RECT 188.675 164.525 189.200 165.050 ;
        RECT 197.175 164.525 197.700 165.050 ;
        RECT 156.650 164.000 197.700 164.525 ;
        RECT 90.725 133.000 91.850 164.000 ;
        RECT 196.350 154.975 197.700 164.000 ;
        RECT 206.200 163.200 207.550 174.025 ;
        RECT 196.350 153.625 207.800 154.975 ;
        RECT 65.000 123.450 201.050 129.375 ;
        RECT 90.145 122.925 90.670 123.450 ;
        RECT 98.645 122.925 99.170 123.450 ;
        RECT 107.120 122.925 107.645 123.450 ;
        RECT 115.620 122.925 116.145 123.450 ;
        RECT 124.095 122.925 124.620 123.450 ;
        RECT 132.595 122.925 133.120 123.450 ;
        RECT 141.070 122.925 141.595 123.450 ;
        RECT 149.570 122.925 150.095 123.450 ;
        RECT 158.045 122.925 158.570 123.450 ;
        RECT 166.545 122.925 167.070 123.450 ;
        RECT 175.045 122.925 175.570 123.450 ;
        RECT 183.520 122.925 184.045 123.450 ;
        RECT 192.020 122.925 192.545 123.450 ;
        RECT 200.520 122.925 201.045 123.450 ;
        RECT 90.140 121.730 90.660 122.925 ;
        RECT 89.095 119.120 91.705 121.730 ;
        RECT 90.140 116.730 90.660 119.120 ;
        RECT 89.095 114.120 91.705 116.730 ;
        RECT 90.140 111.730 90.660 114.120 ;
        RECT 75.275 102.400 81.175 111.300 ;
        RECT 89.095 109.120 91.705 111.730 ;
        RECT 90.140 106.730 90.660 109.120 ;
        RECT 89.095 104.120 91.705 106.730 ;
        RECT 90.140 102.925 90.660 104.120 ;
        RECT 93.340 102.925 93.860 122.925 ;
        RECT 98.630 121.730 99.150 122.925 ;
        RECT 97.585 119.120 100.195 121.730 ;
        RECT 98.630 116.730 99.150 119.120 ;
        RECT 97.585 114.120 100.195 116.730 ;
        RECT 98.630 111.730 99.150 114.120 ;
        RECT 97.585 109.120 100.195 111.730 ;
        RECT 98.630 106.730 99.150 109.120 ;
        RECT 97.585 104.120 100.195 106.730 ;
        RECT 98.630 102.925 99.150 104.120 ;
        RECT 101.830 102.925 102.350 122.925 ;
        RECT 107.120 121.730 107.640 122.925 ;
        RECT 106.075 119.120 108.685 121.730 ;
        RECT 107.120 116.730 107.640 119.120 ;
        RECT 106.075 114.120 108.685 116.730 ;
        RECT 107.120 111.730 107.640 114.120 ;
        RECT 106.075 109.120 108.685 111.730 ;
        RECT 107.120 106.730 107.640 109.120 ;
        RECT 106.075 104.120 108.685 106.730 ;
        RECT 107.120 102.925 107.640 104.120 ;
        RECT 110.320 102.925 110.840 122.925 ;
        RECT 115.610 121.730 116.130 122.925 ;
        RECT 114.565 119.120 117.175 121.730 ;
        RECT 115.610 116.730 116.130 119.120 ;
        RECT 114.565 114.120 117.175 116.730 ;
        RECT 115.610 111.730 116.130 114.120 ;
        RECT 114.565 109.120 117.175 111.730 ;
        RECT 115.610 106.730 116.130 109.120 ;
        RECT 114.565 104.120 117.175 106.730 ;
        RECT 115.610 102.925 116.130 104.120 ;
        RECT 118.810 102.925 119.330 122.925 ;
        RECT 124.100 121.730 124.620 122.925 ;
        RECT 123.055 119.120 125.665 121.730 ;
        RECT 124.100 116.730 124.620 119.120 ;
        RECT 123.055 114.120 125.665 116.730 ;
        RECT 124.100 111.730 124.620 114.120 ;
        RECT 123.055 109.120 125.665 111.730 ;
        RECT 124.100 106.730 124.620 109.120 ;
        RECT 123.055 104.120 125.665 106.730 ;
        RECT 124.100 102.925 124.620 104.120 ;
        RECT 127.300 102.925 127.820 122.925 ;
        RECT 132.590 121.730 133.110 122.925 ;
        RECT 131.545 119.120 134.155 121.730 ;
        RECT 132.590 116.730 133.110 119.120 ;
        RECT 131.545 114.120 134.155 116.730 ;
        RECT 132.590 111.730 133.110 114.120 ;
        RECT 131.545 109.120 134.155 111.730 ;
        RECT 132.590 106.730 133.110 109.120 ;
        RECT 131.545 104.120 134.155 106.730 ;
        RECT 132.590 102.925 133.110 104.120 ;
        RECT 135.790 102.925 136.310 122.925 ;
        RECT 141.080 121.730 141.600 122.925 ;
        RECT 140.035 119.120 142.645 121.730 ;
        RECT 141.080 116.730 141.600 119.120 ;
        RECT 140.035 114.120 142.645 116.730 ;
        RECT 141.080 111.730 141.600 114.120 ;
        RECT 140.035 109.120 142.645 111.730 ;
        RECT 141.080 106.730 141.600 109.120 ;
        RECT 140.035 104.120 142.645 106.730 ;
        RECT 141.080 102.925 141.600 104.120 ;
        RECT 144.280 102.925 144.800 122.925 ;
        RECT 149.570 121.730 150.090 122.925 ;
        RECT 148.525 119.120 151.135 121.730 ;
        RECT 149.570 116.730 150.090 119.120 ;
        RECT 148.525 114.120 151.135 116.730 ;
        RECT 149.570 111.730 150.090 114.120 ;
        RECT 148.525 109.120 151.135 111.730 ;
        RECT 149.570 106.730 150.090 109.120 ;
        RECT 148.525 104.120 151.135 106.730 ;
        RECT 149.570 102.925 150.090 104.120 ;
        RECT 152.770 102.925 153.290 122.925 ;
        RECT 158.060 121.730 158.580 122.925 ;
        RECT 157.015 119.120 159.625 121.730 ;
        RECT 158.060 116.730 158.580 119.120 ;
        RECT 157.015 114.120 159.625 116.730 ;
        RECT 158.060 111.730 158.580 114.120 ;
        RECT 157.015 109.120 159.625 111.730 ;
        RECT 158.060 106.730 158.580 109.120 ;
        RECT 157.015 104.120 159.625 106.730 ;
        RECT 158.060 102.925 158.580 104.120 ;
        RECT 161.260 102.925 161.780 122.925 ;
        RECT 166.550 121.730 167.070 122.925 ;
        RECT 165.505 119.120 168.115 121.730 ;
        RECT 166.550 116.730 167.070 119.120 ;
        RECT 165.505 114.120 168.115 116.730 ;
        RECT 166.550 111.730 167.070 114.120 ;
        RECT 165.505 109.120 168.115 111.730 ;
        RECT 166.550 106.730 167.070 109.120 ;
        RECT 165.505 104.120 168.115 106.730 ;
        RECT 166.550 102.925 167.070 104.120 ;
        RECT 169.750 102.925 170.270 122.925 ;
        RECT 175.040 121.730 175.560 122.925 ;
        RECT 173.995 119.120 176.605 121.730 ;
        RECT 175.040 116.730 175.560 119.120 ;
        RECT 173.995 114.120 176.605 116.730 ;
        RECT 175.040 111.730 175.560 114.120 ;
        RECT 173.995 109.120 176.605 111.730 ;
        RECT 175.040 106.730 175.560 109.120 ;
        RECT 173.995 104.120 176.605 106.730 ;
        RECT 175.040 102.925 175.560 104.120 ;
        RECT 178.240 102.925 178.760 122.925 ;
        RECT 183.530 121.730 184.050 122.925 ;
        RECT 182.485 119.120 185.095 121.730 ;
        RECT 183.530 116.730 184.050 119.120 ;
        RECT 182.485 114.120 185.095 116.730 ;
        RECT 183.530 111.730 184.050 114.120 ;
        RECT 182.485 109.120 185.095 111.730 ;
        RECT 183.530 106.730 184.050 109.120 ;
        RECT 182.485 104.120 185.095 106.730 ;
        RECT 183.530 102.925 184.050 104.120 ;
        RECT 186.730 102.925 187.250 122.925 ;
        RECT 192.020 121.730 192.540 122.925 ;
        RECT 190.975 119.120 193.585 121.730 ;
        RECT 192.020 116.730 192.540 119.120 ;
        RECT 190.975 114.120 193.585 116.730 ;
        RECT 192.020 111.730 192.540 114.120 ;
        RECT 190.975 109.120 193.585 111.730 ;
        RECT 192.020 106.730 192.540 109.120 ;
        RECT 190.975 104.120 193.585 106.730 ;
        RECT 192.020 102.925 192.540 104.120 ;
        RECT 195.220 102.925 195.740 122.925 ;
        RECT 200.510 121.730 201.030 122.925 ;
        RECT 199.465 119.120 202.075 121.730 ;
        RECT 200.510 116.730 201.030 119.120 ;
        RECT 199.465 114.120 202.075 116.730 ;
        RECT 200.510 111.730 201.030 114.120 ;
        RECT 199.465 109.120 202.075 111.730 ;
        RECT 200.510 106.730 201.030 109.120 ;
        RECT 199.465 104.120 202.075 106.730 ;
        RECT 200.510 102.925 201.030 104.120 ;
        RECT 203.710 102.925 204.230 122.925 ;
        RECT 206.450 122.025 207.800 153.625 ;
        RECT 210.000 126.225 211.350 174.675 ;
        RECT 214.625 174.525 215.150 175.050 ;
        RECT 214.600 174.025 215.175 174.525 ;
        RECT 214.125 124.100 215.475 174.025 ;
        RECT 213.850 122.025 215.700 124.100 ;
        RECT 93.345 102.400 93.870 102.925 ;
        RECT 101.820 102.400 102.345 102.925 ;
        RECT 110.320 102.400 110.845 102.925 ;
        RECT 118.820 102.400 119.345 102.925 ;
        RECT 127.295 102.400 127.820 102.925 ;
        RECT 135.795 102.400 136.320 102.925 ;
        RECT 144.270 102.400 144.795 102.925 ;
        RECT 152.770 102.400 153.295 102.925 ;
        RECT 161.270 102.400 161.795 102.925 ;
        RECT 169.745 102.400 170.270 102.925 ;
        RECT 178.245 102.400 178.770 102.925 ;
        RECT 186.720 102.400 187.245 102.925 ;
        RECT 195.220 102.400 195.745 102.925 ;
        RECT 203.695 102.400 204.220 102.925 ;
        RECT 75.275 96.475 204.225 102.400 ;
        RECT 82.400 62.100 83.525 92.600 ;
        RECT 206.450 72.275 207.800 103.825 ;
        RECT 213.975 101.750 215.825 103.825 ;
        RECT 193.150 70.925 207.800 72.275 ;
        RECT 193.150 62.100 194.500 70.925 ;
        RECT 69.435 61.575 144.485 62.100 ;
        RECT 69.435 61.050 69.960 61.575 ;
        RECT 77.935 61.050 78.460 61.575 ;
        RECT 86.410 61.050 86.935 61.575 ;
        RECT 94.910 61.050 95.435 61.575 ;
        RECT 103.385 61.050 103.910 61.575 ;
        RECT 110.010 61.050 110.535 61.575 ;
        RECT 118.485 61.050 119.010 61.575 ;
        RECT 126.985 61.050 127.510 61.575 ;
        RECT 135.460 61.050 135.985 61.575 ;
        RECT 143.960 61.050 144.485 61.575 ;
        RECT 153.450 61.575 194.500 62.100 ;
        RECT 153.450 61.050 153.975 61.575 ;
        RECT 161.950 61.050 162.475 61.575 ;
        RECT 170.425 61.050 170.950 61.575 ;
        RECT 177.000 61.050 177.525 61.575 ;
        RECT 185.475 61.050 186.000 61.575 ;
        RECT 193.975 61.050 194.500 61.575 ;
        RECT 69.440 59.855 69.960 61.050 ;
        RECT 68.395 57.245 71.005 59.855 ;
        RECT 69.440 54.855 69.960 57.245 ;
        RECT 68.395 52.245 71.005 54.855 ;
        RECT 69.440 49.855 69.960 52.245 ;
        RECT 68.395 47.245 71.005 49.855 ;
        RECT 69.440 44.855 69.960 47.245 ;
        RECT 68.395 42.245 71.005 44.855 ;
        RECT 69.440 39.855 69.960 42.245 ;
        RECT 68.395 37.245 71.005 39.855 ;
        RECT 69.440 34.855 69.960 37.245 ;
        RECT 68.395 32.245 71.005 34.855 ;
        RECT 69.440 29.855 69.960 32.245 ;
        RECT 68.395 27.245 71.005 29.855 ;
        RECT 69.440 26.050 69.960 27.245 ;
        RECT 72.640 26.050 73.160 61.050 ;
        RECT 77.930 59.855 78.450 61.050 ;
        RECT 76.885 57.245 79.495 59.855 ;
        RECT 77.930 54.855 78.450 57.245 ;
        RECT 76.885 52.245 79.495 54.855 ;
        RECT 77.930 49.855 78.450 52.245 ;
        RECT 76.885 47.245 79.495 49.855 ;
        RECT 77.930 44.855 78.450 47.245 ;
        RECT 76.885 42.245 79.495 44.855 ;
        RECT 77.930 39.855 78.450 42.245 ;
        RECT 76.885 37.245 79.495 39.855 ;
        RECT 77.930 34.855 78.450 37.245 ;
        RECT 76.885 32.245 79.495 34.855 ;
        RECT 77.930 29.855 78.450 32.245 ;
        RECT 76.885 27.245 79.495 29.855 ;
        RECT 77.930 26.050 78.450 27.245 ;
        RECT 81.130 26.050 81.650 61.050 ;
        RECT 86.420 59.855 86.940 61.050 ;
        RECT 85.375 57.245 87.985 59.855 ;
        RECT 86.420 54.855 86.940 57.245 ;
        RECT 85.375 52.245 87.985 54.855 ;
        RECT 86.420 49.855 86.940 52.245 ;
        RECT 85.375 47.245 87.985 49.855 ;
        RECT 86.420 44.855 86.940 47.245 ;
        RECT 85.375 42.245 87.985 44.855 ;
        RECT 86.420 39.855 86.940 42.245 ;
        RECT 85.375 37.245 87.985 39.855 ;
        RECT 86.420 34.855 86.940 37.245 ;
        RECT 85.375 32.245 87.985 34.855 ;
        RECT 86.420 29.855 86.940 32.245 ;
        RECT 85.375 27.245 87.985 29.855 ;
        RECT 86.420 26.050 86.940 27.245 ;
        RECT 89.620 26.050 90.140 61.050 ;
        RECT 94.910 59.855 95.430 61.050 ;
        RECT 93.865 57.245 96.475 59.855 ;
        RECT 94.910 54.855 95.430 57.245 ;
        RECT 93.865 52.245 96.475 54.855 ;
        RECT 94.910 49.855 95.430 52.245 ;
        RECT 93.865 47.245 96.475 49.855 ;
        RECT 94.910 44.855 95.430 47.245 ;
        RECT 93.865 42.245 96.475 44.855 ;
        RECT 94.910 39.855 95.430 42.245 ;
        RECT 93.865 37.245 96.475 39.855 ;
        RECT 94.910 34.855 95.430 37.245 ;
        RECT 93.865 32.245 96.475 34.855 ;
        RECT 94.910 29.855 95.430 32.245 ;
        RECT 93.865 27.245 96.475 29.855 ;
        RECT 94.910 26.050 95.430 27.245 ;
        RECT 98.110 26.050 98.630 61.050 ;
        RECT 103.400 59.855 103.920 61.050 ;
        RECT 102.355 57.245 104.965 59.855 ;
        RECT 103.400 54.855 103.920 57.245 ;
        RECT 102.355 52.245 104.965 54.855 ;
        RECT 103.400 49.855 103.920 52.245 ;
        RECT 102.355 47.245 104.965 49.855 ;
        RECT 103.400 44.855 103.920 47.245 ;
        RECT 102.355 42.245 104.965 44.855 ;
        RECT 103.400 39.855 103.920 42.245 ;
        RECT 102.355 37.245 104.965 39.855 ;
        RECT 103.400 34.855 103.920 37.245 ;
        RECT 102.355 32.245 104.965 34.855 ;
        RECT 103.400 29.855 103.920 32.245 ;
        RECT 102.355 27.245 104.965 29.855 ;
        RECT 103.400 26.050 103.920 27.245 ;
        RECT 106.600 26.050 107.120 61.050 ;
        RECT 110.000 26.050 110.520 61.050 ;
        RECT 113.200 59.855 113.720 61.050 ;
        RECT 112.155 57.245 114.765 59.855 ;
        RECT 113.200 54.855 113.720 57.245 ;
        RECT 112.155 52.245 114.765 54.855 ;
        RECT 113.200 49.855 113.720 52.245 ;
        RECT 112.155 47.245 114.765 49.855 ;
        RECT 113.200 44.855 113.720 47.245 ;
        RECT 112.155 42.245 114.765 44.855 ;
        RECT 113.200 39.855 113.720 42.245 ;
        RECT 112.155 37.245 114.765 39.855 ;
        RECT 113.200 34.855 113.720 37.245 ;
        RECT 112.155 32.245 114.765 34.855 ;
        RECT 113.200 29.855 113.720 32.245 ;
        RECT 112.155 27.245 114.765 29.855 ;
        RECT 113.200 26.050 113.720 27.245 ;
        RECT 118.490 26.050 119.010 61.050 ;
        RECT 121.690 59.855 122.210 61.050 ;
        RECT 120.645 57.245 123.255 59.855 ;
        RECT 121.690 54.855 122.210 57.245 ;
        RECT 120.645 52.245 123.255 54.855 ;
        RECT 121.690 49.855 122.210 52.245 ;
        RECT 120.645 47.245 123.255 49.855 ;
        RECT 121.690 44.855 122.210 47.245 ;
        RECT 120.645 42.245 123.255 44.855 ;
        RECT 121.690 39.855 122.210 42.245 ;
        RECT 120.645 37.245 123.255 39.855 ;
        RECT 121.690 34.855 122.210 37.245 ;
        RECT 120.645 32.245 123.255 34.855 ;
        RECT 121.690 29.855 122.210 32.245 ;
        RECT 120.645 27.245 123.255 29.855 ;
        RECT 121.690 26.050 122.210 27.245 ;
        RECT 126.980 26.050 127.500 61.050 ;
        RECT 130.180 59.855 130.700 61.050 ;
        RECT 129.135 57.245 131.745 59.855 ;
        RECT 130.180 54.855 130.700 57.245 ;
        RECT 129.135 52.245 131.745 54.855 ;
        RECT 130.180 49.855 130.700 52.245 ;
        RECT 129.135 47.245 131.745 49.855 ;
        RECT 130.180 44.855 130.700 47.245 ;
        RECT 129.135 42.245 131.745 44.855 ;
        RECT 130.180 39.855 130.700 42.245 ;
        RECT 129.135 37.245 131.745 39.855 ;
        RECT 130.180 34.855 130.700 37.245 ;
        RECT 129.135 32.245 131.745 34.855 ;
        RECT 130.180 29.855 130.700 32.245 ;
        RECT 129.135 27.245 131.745 29.855 ;
        RECT 130.180 26.050 130.700 27.245 ;
        RECT 135.470 26.050 135.990 61.050 ;
        RECT 138.670 59.855 139.190 61.050 ;
        RECT 137.625 57.245 140.235 59.855 ;
        RECT 138.670 54.855 139.190 57.245 ;
        RECT 137.625 52.245 140.235 54.855 ;
        RECT 138.670 49.855 139.190 52.245 ;
        RECT 137.625 47.245 140.235 49.855 ;
        RECT 138.670 44.855 139.190 47.245 ;
        RECT 137.625 42.245 140.235 44.855 ;
        RECT 138.670 39.855 139.190 42.245 ;
        RECT 137.625 37.245 140.235 39.855 ;
        RECT 138.670 34.855 139.190 37.245 ;
        RECT 137.625 32.245 140.235 34.855 ;
        RECT 138.670 29.855 139.190 32.245 ;
        RECT 137.625 27.245 140.235 29.855 ;
        RECT 138.670 26.050 139.190 27.245 ;
        RECT 143.960 26.050 144.480 61.050 ;
        RECT 147.160 59.855 147.680 61.050 ;
        RECT 153.440 59.855 153.960 61.050 ;
        RECT 146.115 57.245 148.725 59.855 ;
        RECT 152.395 57.245 155.005 59.855 ;
        RECT 147.160 54.855 147.680 57.245 ;
        RECT 153.440 54.855 153.960 57.245 ;
        RECT 146.115 52.245 148.725 54.855 ;
        RECT 152.395 52.245 155.005 54.855 ;
        RECT 147.160 49.855 147.680 52.245 ;
        RECT 153.440 49.855 153.960 52.245 ;
        RECT 146.115 47.245 148.725 49.855 ;
        RECT 152.395 47.245 155.005 49.855 ;
        RECT 147.160 44.855 147.680 47.245 ;
        RECT 153.440 44.855 153.960 47.245 ;
        RECT 146.115 42.245 148.725 44.855 ;
        RECT 152.395 42.245 155.005 44.855 ;
        RECT 147.160 39.855 147.680 42.245 ;
        RECT 153.440 39.855 153.960 42.245 ;
        RECT 146.115 37.245 148.725 39.855 ;
        RECT 152.395 37.245 155.005 39.855 ;
        RECT 147.160 34.855 147.680 37.245 ;
        RECT 153.440 34.855 153.960 37.245 ;
        RECT 146.115 32.245 148.725 34.855 ;
        RECT 152.395 32.245 155.005 34.855 ;
        RECT 147.160 29.855 147.680 32.245 ;
        RECT 153.440 29.855 153.960 32.245 ;
        RECT 146.115 27.245 148.725 29.855 ;
        RECT 152.395 27.245 155.005 29.855 ;
        RECT 147.160 26.050 147.680 27.245 ;
        RECT 153.440 26.050 153.960 27.245 ;
        RECT 156.640 26.050 157.160 61.050 ;
        RECT 161.930 59.855 162.450 61.050 ;
        RECT 160.885 57.245 163.495 59.855 ;
        RECT 161.930 54.855 162.450 57.245 ;
        RECT 160.885 52.245 163.495 54.855 ;
        RECT 161.930 49.855 162.450 52.245 ;
        RECT 160.885 47.245 163.495 49.855 ;
        RECT 161.930 44.855 162.450 47.245 ;
        RECT 160.885 42.245 163.495 44.855 ;
        RECT 161.930 39.855 162.450 42.245 ;
        RECT 160.885 37.245 163.495 39.855 ;
        RECT 161.930 34.855 162.450 37.245 ;
        RECT 160.885 32.245 163.495 34.855 ;
        RECT 161.930 29.855 162.450 32.245 ;
        RECT 160.885 27.245 163.495 29.855 ;
        RECT 161.930 26.050 162.450 27.245 ;
        RECT 165.130 26.050 165.650 61.050 ;
        RECT 170.420 59.855 170.940 61.050 ;
        RECT 169.375 57.245 171.985 59.855 ;
        RECT 170.420 54.855 170.940 57.245 ;
        RECT 169.375 52.245 171.985 54.855 ;
        RECT 170.420 49.855 170.940 52.245 ;
        RECT 169.375 47.245 171.985 49.855 ;
        RECT 170.420 44.855 170.940 47.245 ;
        RECT 169.375 42.245 171.985 44.855 ;
        RECT 170.420 39.855 170.940 42.245 ;
        RECT 169.375 37.245 171.985 39.855 ;
        RECT 170.420 34.855 170.940 37.245 ;
        RECT 169.375 32.245 171.985 34.855 ;
        RECT 170.420 29.855 170.940 32.245 ;
        RECT 169.375 27.245 171.985 29.855 ;
        RECT 170.420 26.050 170.940 27.245 ;
        RECT 173.620 26.050 174.140 61.050 ;
        RECT 177.010 26.050 177.530 61.050 ;
        RECT 180.210 59.855 180.730 61.050 ;
        RECT 179.165 57.245 181.775 59.855 ;
        RECT 180.210 54.855 180.730 57.245 ;
        RECT 179.165 52.245 181.775 54.855 ;
        RECT 180.210 49.855 180.730 52.245 ;
        RECT 179.165 47.245 181.775 49.855 ;
        RECT 180.210 44.855 180.730 47.245 ;
        RECT 179.165 42.245 181.775 44.855 ;
        RECT 180.210 39.855 180.730 42.245 ;
        RECT 179.165 37.245 181.775 39.855 ;
        RECT 180.210 34.855 180.730 37.245 ;
        RECT 179.165 32.245 181.775 34.855 ;
        RECT 180.210 29.855 180.730 32.245 ;
        RECT 179.165 27.245 181.775 29.855 ;
        RECT 180.210 26.050 180.730 27.245 ;
        RECT 185.500 26.050 186.020 61.050 ;
        RECT 188.700 59.855 189.220 61.050 ;
        RECT 187.655 57.245 190.265 59.855 ;
        RECT 188.700 54.855 189.220 57.245 ;
        RECT 187.655 52.245 190.265 54.855 ;
        RECT 188.700 49.855 189.220 52.245 ;
        RECT 187.655 47.245 190.265 49.855 ;
        RECT 188.700 44.855 189.220 47.245 ;
        RECT 187.655 42.245 190.265 44.855 ;
        RECT 188.700 39.855 189.220 42.245 ;
        RECT 187.655 37.245 190.265 39.855 ;
        RECT 188.700 34.855 189.220 37.245 ;
        RECT 187.655 32.245 190.265 34.855 ;
        RECT 188.700 29.855 189.220 32.245 ;
        RECT 187.655 27.245 190.265 29.855 ;
        RECT 188.700 26.050 189.220 27.245 ;
        RECT 193.990 26.050 194.510 61.050 ;
        RECT 197.190 59.855 197.710 61.050 ;
        RECT 196.145 57.245 198.755 59.855 ;
        RECT 197.190 54.855 197.710 57.245 ;
        RECT 196.145 52.245 198.755 54.855 ;
        RECT 203.125 52.550 204.250 53.275 ;
        RECT 197.190 49.855 197.710 52.245 ;
        RECT 203.400 51.575 203.975 52.550 ;
        RECT 203.425 51.050 203.950 51.575 ;
        RECT 203.440 49.855 203.960 51.050 ;
        RECT 206.225 50.825 207.575 62.575 ;
        RECT 210.000 52.725 211.350 99.650 ;
        RECT 210.000 52.100 211.975 52.725 ;
        RECT 211.400 51.575 211.975 52.100 ;
        RECT 211.425 51.050 211.950 51.575 ;
        RECT 196.145 47.245 198.755 49.855 ;
        RECT 202.395 47.245 205.005 49.855 ;
        RECT 197.190 44.855 197.710 47.245 ;
        RECT 203.440 44.855 203.960 47.245 ;
        RECT 196.145 42.245 198.755 44.855 ;
        RECT 202.395 42.245 205.005 44.855 ;
        RECT 197.190 39.855 197.710 42.245 ;
        RECT 203.440 39.855 203.960 42.245 ;
        RECT 196.145 37.245 198.755 39.855 ;
        RECT 202.395 37.245 205.005 39.855 ;
        RECT 197.190 34.855 197.710 37.245 ;
        RECT 203.440 34.855 203.960 37.245 ;
        RECT 196.145 32.245 198.755 34.855 ;
        RECT 202.395 32.245 205.005 34.855 ;
        RECT 197.190 29.855 197.710 32.245 ;
        RECT 203.440 29.855 203.960 32.245 ;
        RECT 196.145 27.245 198.755 29.855 ;
        RECT 202.395 27.245 205.005 29.855 ;
        RECT 197.190 26.050 197.710 27.245 ;
        RECT 203.440 26.050 203.960 27.245 ;
        RECT 206.640 26.050 207.160 50.825 ;
        RECT 211.440 49.855 211.960 51.050 ;
        RECT 214.225 50.950 215.575 101.750 ;
        RECT 210.395 47.245 213.005 49.855 ;
        RECT 211.440 44.855 211.960 47.245 ;
        RECT 210.395 42.245 213.005 44.855 ;
        RECT 211.440 39.855 211.960 42.245 ;
        RECT 210.395 37.245 213.005 39.855 ;
        RECT 211.440 34.855 211.960 37.245 ;
        RECT 210.395 32.245 213.005 34.855 ;
        RECT 211.440 29.855 211.960 32.245 ;
        RECT 210.395 27.245 213.005 29.855 ;
        RECT 211.440 26.050 211.960 27.245 ;
        RECT 214.640 26.050 215.160 50.950 ;
        RECT 72.635 25.525 73.160 26.050 ;
        RECT 81.135 25.525 81.660 26.050 ;
        RECT 89.610 25.525 90.135 26.050 ;
        RECT 98.110 25.525 98.635 26.050 ;
        RECT 106.585 25.525 107.110 26.050 ;
        RECT 113.210 25.525 113.735 26.050 ;
        RECT 121.685 25.525 122.210 26.050 ;
        RECT 130.185 25.525 130.710 26.050 ;
        RECT 138.660 25.525 139.185 26.050 ;
        RECT 147.160 25.525 147.685 26.050 ;
        RECT 72.635 25.000 147.685 25.525 ;
        RECT 156.650 25.525 157.175 26.050 ;
        RECT 165.150 25.525 165.675 26.050 ;
        RECT 173.625 25.525 174.150 26.050 ;
        RECT 180.200 25.525 180.725 26.050 ;
        RECT 188.675 25.525 189.200 26.050 ;
        RECT 197.175 25.525 197.700 26.050 ;
        RECT 206.625 25.525 207.150 26.050 ;
        RECT 214.625 25.525 215.150 26.050 ;
        RECT 156.650 25.000 197.700 25.525 ;
        RECT 206.600 25.000 207.175 25.525 ;
        RECT 214.600 25.000 215.175 25.525 ;
        RECT 73.400 5.650 75.425 7.575 ;
        RECT 92.725 5.650 94.750 12.775 ;
        RECT 112.050 5.650 114.075 18.125 ;
        RECT 131.375 5.650 133.400 23.400 ;
        RECT 74.525 1.000 75.425 5.650 ;
        RECT 93.850 1.000 94.750 5.650 ;
        RECT 113.150 1.000 114.075 5.650 ;
        RECT 132.475 1.000 133.400 5.650 ;
        RECT 151.800 5.650 154.775 8.700 ;
        RECT 151.800 1.000 152.725 5.650 ;
  END
END tt_um_TinyWhisper
END LIBRARY

