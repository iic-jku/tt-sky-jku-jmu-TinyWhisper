magic
tech sky130A
magscale 1 2
timestamp 1762641840
<< locali >>
rect -5115 5305 25055 5770
rect -3235 3170 -2950 5305
rect -575 3170 -290 5305
rect 2060 3170 2440 5305
rect 4220 3170 4550 5305
rect 6880 3170 7210 5305
rect 9555 3170 9885 5305
rect 12215 3170 12545 5305
rect 14865 3170 15195 5305
rect 17555 3170 17885 5305
rect 19690 3170 20020 5305
rect 22340 3170 22670 5305
rect -3250 2145 -2925 3060
rect -640 2145 -225 3060
rect 2090 2145 2405 3060
rect 4205 2145 4535 3060
rect 6900 2145 7205 3060
rect 9575 2145 9895 3060
rect 12220 2145 12585 3060
rect 14755 2145 15330 3060
rect 17420 2145 17990 3060
rect 19570 2145 20145 3060
rect 22235 2145 22810 3060
rect -5115 1680 25055 2145
<< metal1 >>
rect -5165 5620 25055 5770
rect -3035 3260 -2840 3270
rect -5165 3060 -5115 3170
rect -3035 2970 -3025 3260
rect -2850 2970 -2840 3260
rect -3035 2960 -2840 2970
rect -370 3260 -100 3270
rect -370 2970 -360 3260
rect -185 2970 -100 3260
rect -370 2960 -100 2970
rect 1980 3260 2565 3270
rect 1980 2970 1990 3260
rect 2480 2970 2565 3260
rect 3795 3160 3990 3300
rect 3980 3070 3990 3160
rect 3040 3065 3780 3070
rect 1980 2960 2565 2970
rect 3795 2925 3990 3070
rect 4445 3260 4715 3270
rect 4445 2970 4455 3260
rect 4630 2970 4715 3260
rect 4445 2960 4715 2970
rect 7110 3260 7380 3270
rect 7110 2970 7120 3260
rect 7295 2970 7380 3260
rect 7110 2960 7380 2970
rect 9775 3260 10045 3270
rect 9775 2970 9785 3260
rect 9960 2970 10045 3260
rect 9775 2960 10045 2970
rect 12440 3260 12710 3270
rect 12440 2970 12450 3260
rect 12625 2970 12710 3260
rect 12440 2960 12710 2970
rect 15105 3260 15375 3270
rect 15105 2970 15115 3260
rect 15290 2970 15375 3260
rect 15105 2960 15375 2970
rect 17770 3260 18040 3270
rect 17770 2970 17780 3260
rect 17955 2970 18040 3260
rect 18515 3065 19255 3070
rect 17770 2960 18040 2970
rect 19265 2925 19465 3305
rect 19920 3260 20190 3270
rect 19920 2970 19930 3260
rect 20105 2970 20190 3260
rect 19920 2960 20190 2970
rect 22585 3260 22855 3270
rect 22585 2970 22595 3260
rect 22770 2970 22855 3260
rect 22585 2960 22855 2970
rect -5165 1680 25055 1830
<< via1 >>
rect -3025 2970 -2850 3260
rect -360 2970 -185 3260
rect 1990 2970 2480 3260
rect 2980 3070 3980 3160
rect 4455 2970 4630 3260
rect 7120 2970 7295 3260
rect 9785 2970 9960 3260
rect 12450 2970 12625 3260
rect 15115 2970 15290 3260
rect 17780 2970 17955 3260
rect 18515 3070 19255 3130
rect 19930 2970 20105 3260
rect 22595 2970 22770 3260
<< metal2 >>
rect -3305 5375 24850 5525
rect -3305 2915 -3155 5375
rect -800 4455 -300 4465
rect -800 4165 -555 4455
rect -310 4165 -300 4455
rect -800 4155 -300 4165
rect 1865 4455 2365 4465
rect 1865 4165 2110 4455
rect 2355 4165 2365 4455
rect 1865 4155 2365 4165
rect 6675 4455 7180 4465
rect 6675 4165 6925 4455
rect 7170 4165 7180 4455
rect 6675 4155 7180 4165
rect 12005 4455 12510 4465
rect 12005 4165 12250 4455
rect 12500 4165 12510 4455
rect 12005 4155 12510 4165
rect 22150 4455 22655 4465
rect 22150 4165 22400 4455
rect 22645 4165 22655 4455
rect 22150 4155 22655 4165
rect 24805 4455 25320 4465
rect 24805 4165 25065 4455
rect 25310 4165 25320 4455
rect 24805 4155 25320 4165
rect -3035 3260 -2840 3270
rect -3035 2970 -3025 3260
rect -2850 2970 -2840 3260
rect -3035 2960 -2840 2970
rect -800 2915 -490 4155
rect 1865 3270 2175 4155
rect -370 3260 -175 3270
rect -370 2970 -360 3260
rect -185 2970 -175 3260
rect -370 2960 -175 2970
rect 1865 3260 2490 3270
rect 1865 2970 1990 3260
rect 2480 2970 2490 3260
rect 1865 2960 2490 2970
rect 1865 2915 2175 2960
rect 4010 2720 4320 3315
rect 4445 3260 4640 3270
rect 4445 2970 4455 3260
rect 4630 2970 4640 3260
rect 4445 2960 4640 2970
rect 6675 2915 6985 4155
rect 7110 3260 7305 3270
rect 7110 2970 7120 3260
rect 7295 2970 7305 3260
rect 7110 2960 7305 2970
rect 9340 2720 9650 3315
rect 9775 3260 9970 3270
rect 9775 2970 9785 3260
rect 9960 2970 9970 3260
rect 9775 2960 9970 2970
rect 12005 2915 12315 4155
rect 17335 3745 17840 3755
rect 17335 3455 17585 3745
rect 17830 3455 17840 3745
rect 17335 3445 17840 3455
rect 12440 3260 12635 3270
rect 12440 2970 12450 3260
rect 12625 2970 12635 3260
rect 12440 2960 12635 2970
rect 14670 3260 14980 3315
rect 14670 2970 14680 3260
rect 14970 2970 14980 3260
rect 14670 2915 14980 2970
rect 15105 3260 15300 3270
rect 15105 2970 15115 3260
rect 15290 2970 15300 3260
rect 15105 2960 15300 2970
rect 17335 2915 17645 3445
rect 17770 3260 17965 3270
rect 17770 2970 17780 3260
rect 17955 2970 17965 3260
rect 19920 3260 20115 3270
rect 18455 3130 19455 3160
rect 18455 3070 18515 3130
rect 19255 3070 19455 3130
rect 17770 2960 17965 2970
rect 19920 2970 19930 3260
rect 20105 2970 20115 3260
rect 19920 2960 20115 2970
rect 22150 3260 22460 4155
rect 22150 2970 22160 3260
rect 22450 2970 22460 3260
rect 22150 2915 22460 2970
rect 22585 3260 22780 3270
rect 22585 2970 22595 3260
rect 22770 2970 22780 3260
rect 22585 2960 22780 2970
rect 24805 2915 25115 4155
rect 4010 2710 4515 2720
rect 4010 2420 4260 2710
rect 4505 2420 4515 2710
rect 4010 2410 4515 2420
rect 9340 2710 9845 2720
rect 9340 2420 9590 2710
rect 9835 2420 9845 2710
rect 9340 2410 9845 2420
<< via2 >>
rect -555 4165 -310 4455
rect 2110 4165 2355 4455
rect 6925 4165 7170 4455
rect 12250 4165 12500 4455
rect 22400 4165 22645 4455
rect 25065 4165 25310 4455
rect -3025 2970 -2850 3260
rect -360 2970 -185 3260
rect 4455 2970 4630 3260
rect 7120 2970 7295 3260
rect 9785 2970 9960 3260
rect 17585 3455 17830 3745
rect 12450 2970 12625 3260
rect 14680 2970 14970 3260
rect 15115 2970 15290 3260
rect 17780 2970 17955 3260
rect 19930 2970 20105 3260
rect 22160 2970 22450 3260
rect 22595 2970 22770 3260
rect 4260 2420 4505 2710
rect 9590 2420 9835 2710
<< metal3 >>
rect -3250 5525 4640 5935
rect -3250 3260 -2840 5525
rect -565 4455 2365 4465
rect -565 4165 -555 4455
rect -310 4165 2110 4455
rect 2355 4165 2365 4455
rect -565 4155 2365 4165
rect -3250 2970 -3025 3260
rect -2850 2970 -2840 3260
rect -3250 2960 -2840 2970
rect -585 3260 -175 3270
rect -585 2970 -360 3260
rect -185 2970 -175 3260
rect -585 1925 -175 2970
rect 4230 3260 4640 5525
rect 6895 5525 22995 5935
rect 6895 4455 7205 5525
rect 6895 4165 6925 4455
rect 7170 4165 7205 4455
rect 6895 4155 7205 4165
rect 12225 4455 12535 5525
rect 12225 4165 12250 4455
rect 12500 4165 12535 4455
rect 12225 4155 12535 4165
rect 4230 2970 4455 3260
rect 4630 2970 4640 3260
rect 4230 2960 4640 2970
rect 5550 3745 17840 3755
rect 5550 3455 17585 3745
rect 17830 3455 17840 3745
rect 5550 3445 17840 3455
rect 5550 2720 5860 3445
rect 4250 2710 5860 2720
rect 4250 2420 4260 2710
rect 4505 2420 5860 2710
rect 4250 2410 5860 2420
rect 6895 3260 7305 3270
rect 6895 2970 7120 3260
rect 7295 2970 7305 3260
rect 6895 1925 7305 2970
rect 9560 3260 9970 3445
rect 9560 2970 9785 3260
rect 9960 2970 9970 3260
rect 9560 2960 9970 2970
rect 12225 3260 12635 3445
rect 12225 2970 12450 3260
rect 12625 2970 12635 3260
rect 12225 2960 12635 2970
rect 14570 3260 14980 3315
rect 14570 2970 14680 3260
rect 14970 2970 14980 3260
rect -585 1515 7305 1925
rect 9560 2710 9870 2720
rect 9560 2420 9590 2710
rect 9835 2420 9870 2710
rect 9560 1925 9870 2420
rect 14570 1925 14980 2970
rect 15105 3260 15515 3270
rect 15105 2970 15115 3260
rect 15290 2970 15515 3260
rect 15105 2855 15515 2970
rect 17770 3260 18180 3270
rect 17770 2970 17780 3260
rect 17955 2970 18180 3260
rect 17770 2855 18180 2970
rect 19705 3260 20115 5525
rect 22390 4455 25320 4465
rect 22390 4165 22400 4455
rect 22645 4165 25065 4455
rect 25310 4165 25320 4455
rect 22390 4155 25320 4165
rect 19705 2970 19930 3260
rect 20105 2970 20115 3260
rect 19705 2960 20115 2970
rect 21030 3260 22460 3270
rect 21030 2970 22160 3260
rect 22450 2970 22460 3260
rect 21030 2960 22460 2970
rect 22585 3260 22995 3270
rect 22585 2970 22595 3260
rect 22770 2970 22995 3260
rect 21030 2855 21340 2960
rect 15105 2545 21340 2855
rect 22585 1925 22995 2970
rect 9560 1515 22995 1925
use inverter_lv_en_NF4  inverter_lv_en_NF4_0 inverter/inverter_lv_en_NF4
timestamp 1762641840
transform 1 0 2495 0 1 1075
box -165 605 1770 4695
use inverter_lv_en_NF4  inverter_lv_en_NF4_1
timestamp 1762641840
transform 1 0 17970 0 1 1075
box -165 605 1770 4695
use inverter_lv_en_NF6  inverter_lv_en_NF6_0 inverter/inverter_lv_en_NF6
timestamp 1762641840
transform 1 0 -2835 0 1 1075
box -165 605 2305 4695
use inverter_lv_en_NF6  inverter_lv_en_NF6_1
timestamp 1762641840
transform 1 0 -170 0 1 1075
box -165 605 2305 4695
use inverter_lv_en_NF6  inverter_lv_en_NF6_2
timestamp 1762641840
transform 1 0 4645 0 1 1075
box -165 605 2305 4695
use inverter_lv_en_NF6  inverter_lv_en_NF6_3
timestamp 1762641840
transform 1 0 7310 0 1 1075
box -165 605 2305 4695
use inverter_lv_en_NF6  inverter_lv_en_NF6_4
timestamp 1762641840
transform 1 0 9975 0 1 1075
box -165 605 2305 4695
use inverter_lv_en_NF6  inverter_lv_en_NF6_5
timestamp 1762641840
transform 1 0 12640 0 1 1075
box -165 605 2305 4695
use inverter_lv_en_NF6  inverter_lv_en_NF6_6
timestamp 1762641840
transform 1 0 15305 0 1 1075
box -165 605 2305 4695
use inverter_lv_en_NF6  inverter_lv_en_NF6_7
timestamp 1762641840
transform 1 0 20120 0 1 1075
box -165 605 2305 4695
use inverter_lv_en_NF6  inverter_lv_en_NF6_8
timestamp 1762641840
transform 1 0 22785 0 1 1075
box -165 605 2305 4695
use inverter_lv_NF4  inverter_lv_NF4_0 inverter/inverter_lv_NF4
timestamp 1762641840
transform 1 0 -4985 0 1 1075
box -165 605 1770 4695
<< labels >>
flabel metal1 -5145 1750 -5145 1750 0 FreeSans 400 0 0 0 VSS
port 3 nsew
flabel metal2 -2925 5445 -2925 5445 0 FreeSans 320 0 0 0 ota_core_en_n
flabel metal1 -5155 3110 -5155 3110 0 FreeSans 320 0 0 0 di_ota_core_en
port 20 nsew
flabel metal1 -5150 5695 -5150 5695 0 FreeSans 400 0 0 0 VDD
port 5 nsew
flabel metal3 -2965 5760 -2965 5760 0 FreeSans 1600 0 0 0 vinp
port 30 nsew
flabel metal3 -325 1720 -325 1720 0 FreeSans 1600 0 0 0 vinn
port 32 nsew
flabel metal3 22480 1710 22480 1710 0 FreeSans 1600 0 0 0 voutp
port 40 nsew
flabel metal3 22450 5725 22450 5725 0 FreeSans 1600 0 0 0 voutn
port 42 nsew
<< end >>
