magic
tech sky130A
magscale 1 2
timestamp 1762641840
<< locali >>
rect -2055 6685 2285 7530
rect 25355 6685 28500 7530
rect -2055 6000 2280 6685
rect 26015 6005 28500 6685
rect 28250 2985 28500 6005
rect 28115 1775 28500 2985
rect -2055 965 2280 1645
rect 26015 965 28500 1775
rect -2055 120 2295 965
rect 25420 120 28500 965
<< metal1 >>
rect -2055 7520 2350 7530
rect -2055 7205 -2045 7520
rect -885 7205 2350 7520
rect -2055 6685 2350 7205
rect 8430 6945 8650 7350
rect 25420 6685 28500 7530
rect -2105 6145 2510 6550
rect 5275 6145 5500 6550
rect 25420 6530 25715 6550
rect 25420 6165 25470 6530
rect 25695 6165 25715 6530
rect 25420 6145 25715 6165
rect 26015 6005 28500 6685
rect -2105 5855 -1930 5865
rect -2105 5725 -2045 5855
rect -2105 5715 -1930 5725
rect -2105 5520 -1985 5715
rect -2105 3155 -2055 3265
rect 28250 2985 28500 6005
rect -2055 2390 -1970 2970
rect -2105 2100 -1885 2110
rect -2105 1785 -2045 2100
rect 28115 1805 28500 2985
rect -2105 1775 -1885 1785
rect -2110 1100 2510 1505
rect 5280 1100 5495 1505
rect 18870 1145 18880 1460
rect 25450 1485 25715 1505
rect 18950 1145 18960 1460
rect 25450 1120 25470 1485
rect 25695 1120 25715 1485
rect 25450 1100 25715 1120
rect 26015 965 28500 1805
rect -2055 445 2350 965
rect -2055 130 -2045 445
rect -885 130 2350 445
rect 8430 300 8650 705
rect -2055 120 2350 130
rect 25425 120 28500 965
<< via1 >>
rect -2045 7205 -885 7520
rect 18880 6150 18950 6550
rect 25470 6165 25695 6530
rect -2045 5725 -180 5855
rect 105 5725 2490 5855
rect 2770 5725 5150 5855
rect 5435 5725 7300 5855
rect 7585 5725 9965 5855
rect 10250 5725 12630 5855
rect 12915 5725 15295 5855
rect 15580 5725 17960 5855
rect 18245 5725 20625 5855
rect 20910 5725 22775 5855
rect 23060 5725 25440 5855
rect 25725 5725 28105 5855
rect -2045 1785 -885 2100
rect 18880 1100 18950 1505
rect 25470 1120 25695 1485
rect -2045 130 -885 445
<< metal2 >>
rect -2055 7520 -875 7530
rect -2055 7205 -2045 7520
rect -885 7205 -875 7520
rect -2055 7195 -875 7205
rect 18870 6550 18960 6560
rect 18870 6150 18880 6550
rect 18950 6150 18960 6550
rect 18870 6135 18960 6150
rect 25450 6530 25715 6550
rect 25450 6165 25470 6530
rect 25695 6165 25715 6530
rect 25450 6145 25715 6165
rect -2105 5855 28115 6005
rect -2105 5725 -2045 5855
rect -180 5725 105 5855
rect 2490 5725 2770 5855
rect 5150 5725 5435 5855
rect 7300 5725 7585 5855
rect 9965 5725 10250 5855
rect 12630 5725 12915 5855
rect 15295 5725 15580 5855
rect 17960 5725 18245 5855
rect 20625 5725 20910 5855
rect 22775 5725 23060 5855
rect 25440 5725 25725 5855
rect 28105 5725 28115 5855
rect -2105 5715 28115 5725
rect -2055 2100 -875 2110
rect -2055 1785 -2045 2100
rect -885 1785 -875 2100
rect -2055 1775 -875 1785
rect 18870 1505 18960 1515
rect 18870 1100 18880 1505
rect 18950 1100 18960 1505
rect 25450 1485 25715 1505
rect 25450 1120 25470 1485
rect 25695 1120 25715 1485
rect 25450 1100 25715 1120
rect 18870 1090 18960 1100
rect -2055 445 -875 455
rect -2055 130 -2045 445
rect -885 130 -875 445
rect -2055 120 -875 130
<< via2 >>
rect -2045 7205 -885 7520
rect 18880 6180 18950 6505
rect 25470 6165 25695 6530
rect -2045 1785 -885 2100
rect 18880 1140 18950 1465
rect 25470 1120 25695 1485
rect -2045 130 -885 445
<< metal3 >>
rect -2055 7520 -875 7530
rect -2055 7205 -2045 7520
rect -885 7205 -875 7520
rect -2055 2100 -875 7205
rect 25450 6530 26055 7435
rect 7290 6505 18960 6515
rect 7290 6180 18880 6505
rect 18950 6180 18960 6505
rect 7290 6170 18960 6180
rect 7290 5620 7700 6170
rect 25450 6165 25470 6530
rect 25695 6165 26055 6530
rect 25450 5620 26055 6165
rect -2055 1785 -2045 2100
rect -885 1785 -875 2100
rect -2055 445 -875 1785
rect 9955 1475 10365 1615
rect 25450 1485 26055 2020
rect 9955 1465 18960 1475
rect 9955 1140 18880 1465
rect 18950 1140 18960 1465
rect 9955 1130 18960 1140
rect -2055 130 -2045 445
rect -885 130 -875 445
rect -2055 120 -875 130
rect 25450 1120 25470 1485
rect 25695 1120 26055 1485
rect 25450 120 26055 1120
use ota_core_hybrid_bm  ota_core_hybrid_bm_0 ota_core
timestamp 1762641840
transform 1 0 3061 0 1 94
box -5165 1515 25320 5935
use resistors  resistors_0 resistors
timestamp 1762641840
transform 1 0 2310 0 1 -1385
box -65 1505 23150 8915
<< labels >>
flabel metal1 -1916 1306 -1916 1306 0 FreeSans 1200 0 0 0 vinn
port 5 nsew
flabel metal1 5385 6360 5385 6360 0 FreeSans 400 0 0 0 vC1p
port 29 nsew
flabel metal1 5380 1305 5380 1305 0 FreeSans 400 0 0 0 vC1n
port 31 nsew
flabel metal1 8530 590 8530 590 0 FreeSans 400 0 0 0 vC2n
port 33 nsew
flabel metal1 8540 7150 8540 7150 0 FreeSans 400 0 0 0 vC2p
port 35 nsew
flabel metal1 -2080 3205 -2080 3205 0 FreeSans 400 0 0 0 di_filter_ota_en
port 37 nsew
flabel metal1 -1914 6358 -1914 6358 0 FreeSans 1200 0 0 0 vinp
port 3 nsew
flabel metal1 -2080 5695 -2080 5695 0 FreeSans 1600 0 0 0 VDD
port 52 nsew
flabel metal1 -2080 1955 -2080 1955 0 FreeSans 1600 0 0 0 VSS
port 54 nsew
flabel metal3 25725 405 25725 405 0 FreeSans 1600 0 0 0 voutp
port 58 nsew
flabel metal3 25750 7165 25750 7165 0 FreeSans 1600 0 0 0 voutn
port 60 nsew
<< end >>
