magic
tech sky130A
magscale 1 2
timestamp 1762793988
<< locali >>
rect -33145 12205 -2590 12535
rect -2595 10655 -1985 11275
rect -2595 8625 -1985 9415
rect -2595 6485 -1985 7105
rect -2590 4800 -1980 5245
rect -33145 4455 -1980 4800
<< viali >>
rect -33130 11890 -31980 12195
rect -33130 4815 -31980 5120
<< metal1 >>
rect -33145 12210 -2590 12535
rect -31015 10825 -30480 11230
rect -31940 10220 -31280 10495
rect -2200 10335 -2080 10475
rect -2595 8865 -1975 9205
rect -2595 8860 -1965 8865
rect -2590 8625 -1965 8860
rect -33280 7765 -33175 8015
rect -31790 6470 -31275 6875
rect -30930 5780 -30415 6185
rect -2200 6100 -2080 6290
rect -2595 4800 -1975 5035
rect -33145 4695 -1975 4800
rect -33145 4455 -1970 4695
<< metal2 >>
rect -4920 12265 4565 12535
rect -4920 10405 -3435 12265
<< metal3 >>
rect -5640 12815 3610 13420
rect -5640 12110 -5035 12815
rect 2790 12585 3610 12815
rect 5655 8235 6805 8650
rect -5640 4175 -5035 4815
rect 2790 4175 3610 4405
rect -5640 3565 3610 4175
use passive_voltage_mode_mixer  passive_voltage_mode_mixer_0 passive_voltage_mode_mixer
timestamp 1762641840
transform 1 0 -2200 0 1 8595
box 0 -4195 9030 3995
use third_order_mfb_lp_filter_wo_C  third_order_mfb_lp_filter_wo_C_0 third_order_mfb_lp_filter
timestamp 1762641840
transform 1 0 -31090 0 1 4680
box -2110 120 28500 7530
<< labels >>
flabel metal3 6240 8485 6240 8485 0 FreeSans 1600 0 0 0 vout_RF
port 15 nsew
flabel metal1 -30680 5980 -30680 5980 0 FreeSans 1600 0 0 0 vinn
port 62 nsew
flabel metal1 -30745 11025 -30745 11025 0 FreeSans 1600 0 0 0 vinp
port 68 nsew
flabel metal1 -2145 6215 -2145 6215 0 FreeSans 800 0 0 0 vinp_LO
port 72 nsew
flabel metal1 -2140 10420 -2140 10420 0 FreeSans 800 0 0 0 vinn_LO
port 74 nsew
flabel metal1 -31610 10350 -31610 10350 0 FreeSans 1600 0 0 0 VDD
port 112 nsew
flabel metal1 -33235 7885 -33235 7885 0 FreeSans 1600 0 0 0 di_afe_en
port 114 nsew
flabel metal1 -31645 6635 -31645 6635 0 FreeSans 1600 0 0 0 VSS
port 118 nsew
<< end >>
