magic
tech sky130A
magscale 1 2
timestamp 1762792518
<< nwell >>
rect -2696 -21045 2696 21045
<< pmos >>
rect -2500 15826 2500 20826
rect -2500 10590 2500 15590
rect -2500 5354 2500 10354
rect -2500 118 2500 5118
rect -2500 -5118 2500 -118
rect -2500 -10354 2500 -5354
rect -2500 -15590 2500 -10590
rect -2500 -20826 2500 -15826
<< pdiff >>
rect -2558 20814 -2500 20826
rect -2558 15838 -2546 20814
rect -2512 15838 -2500 20814
rect -2558 15826 -2500 15838
rect 2500 20814 2558 20826
rect 2500 15838 2512 20814
rect 2546 15838 2558 20814
rect 2500 15826 2558 15838
rect -2558 15578 -2500 15590
rect -2558 10602 -2546 15578
rect -2512 10602 -2500 15578
rect -2558 10590 -2500 10602
rect 2500 15578 2558 15590
rect 2500 10602 2512 15578
rect 2546 10602 2558 15578
rect 2500 10590 2558 10602
rect -2558 10342 -2500 10354
rect -2558 5366 -2546 10342
rect -2512 5366 -2500 10342
rect -2558 5354 -2500 5366
rect 2500 10342 2558 10354
rect 2500 5366 2512 10342
rect 2546 5366 2558 10342
rect 2500 5354 2558 5366
rect -2558 5106 -2500 5118
rect -2558 130 -2546 5106
rect -2512 130 -2500 5106
rect -2558 118 -2500 130
rect 2500 5106 2558 5118
rect 2500 130 2512 5106
rect 2546 130 2558 5106
rect 2500 118 2558 130
rect -2558 -130 -2500 -118
rect -2558 -5106 -2546 -130
rect -2512 -5106 -2500 -130
rect -2558 -5118 -2500 -5106
rect 2500 -130 2558 -118
rect 2500 -5106 2512 -130
rect 2546 -5106 2558 -130
rect 2500 -5118 2558 -5106
rect -2558 -5366 -2500 -5354
rect -2558 -10342 -2546 -5366
rect -2512 -10342 -2500 -5366
rect -2558 -10354 -2500 -10342
rect 2500 -5366 2558 -5354
rect 2500 -10342 2512 -5366
rect 2546 -10342 2558 -5366
rect 2500 -10354 2558 -10342
rect -2558 -10602 -2500 -10590
rect -2558 -15578 -2546 -10602
rect -2512 -15578 -2500 -10602
rect -2558 -15590 -2500 -15578
rect 2500 -10602 2558 -10590
rect 2500 -15578 2512 -10602
rect 2546 -15578 2558 -10602
rect 2500 -15590 2558 -15578
rect -2558 -15838 -2500 -15826
rect -2558 -20814 -2546 -15838
rect -2512 -20814 -2500 -15838
rect -2558 -20826 -2500 -20814
rect 2500 -15838 2558 -15826
rect 2500 -20814 2512 -15838
rect 2546 -20814 2558 -15838
rect 2500 -20826 2558 -20814
<< pdiffc >>
rect -2546 15838 -2512 20814
rect 2512 15838 2546 20814
rect -2546 10602 -2512 15578
rect 2512 10602 2546 15578
rect -2546 5366 -2512 10342
rect 2512 5366 2546 10342
rect -2546 130 -2512 5106
rect 2512 130 2546 5106
rect -2546 -5106 -2512 -130
rect 2512 -5106 2546 -130
rect -2546 -10342 -2512 -5366
rect 2512 -10342 2546 -5366
rect -2546 -15578 -2512 -10602
rect 2512 -15578 2546 -10602
rect -2546 -20814 -2512 -15838
rect 2512 -20814 2546 -15838
<< nsubdiff >>
rect -2660 20975 -2564 21009
rect 2564 20975 2660 21009
rect -2660 20913 -2626 20975
rect 2626 20913 2660 20975
rect -2660 -20975 -2626 -20913
rect 2626 -20975 2660 -20913
rect -2660 -21009 -2564 -20975
rect 2564 -21009 2660 -20975
<< nsubdiffcont >>
rect -2564 20975 2564 21009
rect -2660 -20913 -2626 20913
rect 2626 -20913 2660 20913
rect -2564 -21009 2564 -20975
<< poly >>
rect -2500 20907 2500 20923
rect -2500 20873 -2484 20907
rect 2484 20873 2500 20907
rect -2500 20826 2500 20873
rect -2500 15779 2500 15826
rect -2500 15745 -2484 15779
rect 2484 15745 2500 15779
rect -2500 15729 2500 15745
rect -2500 15671 2500 15687
rect -2500 15637 -2484 15671
rect 2484 15637 2500 15671
rect -2500 15590 2500 15637
rect -2500 10543 2500 10590
rect -2500 10509 -2484 10543
rect 2484 10509 2500 10543
rect -2500 10493 2500 10509
rect -2500 10435 2500 10451
rect -2500 10401 -2484 10435
rect 2484 10401 2500 10435
rect -2500 10354 2500 10401
rect -2500 5307 2500 5354
rect -2500 5273 -2484 5307
rect 2484 5273 2500 5307
rect -2500 5257 2500 5273
rect -2500 5199 2500 5215
rect -2500 5165 -2484 5199
rect 2484 5165 2500 5199
rect -2500 5118 2500 5165
rect -2500 71 2500 118
rect -2500 37 -2484 71
rect 2484 37 2500 71
rect -2500 21 2500 37
rect -2500 -37 2500 -21
rect -2500 -71 -2484 -37
rect 2484 -71 2500 -37
rect -2500 -118 2500 -71
rect -2500 -5165 2500 -5118
rect -2500 -5199 -2484 -5165
rect 2484 -5199 2500 -5165
rect -2500 -5215 2500 -5199
rect -2500 -5273 2500 -5257
rect -2500 -5307 -2484 -5273
rect 2484 -5307 2500 -5273
rect -2500 -5354 2500 -5307
rect -2500 -10401 2500 -10354
rect -2500 -10435 -2484 -10401
rect 2484 -10435 2500 -10401
rect -2500 -10451 2500 -10435
rect -2500 -10509 2500 -10493
rect -2500 -10543 -2484 -10509
rect 2484 -10543 2500 -10509
rect -2500 -10590 2500 -10543
rect -2500 -15637 2500 -15590
rect -2500 -15671 -2484 -15637
rect 2484 -15671 2500 -15637
rect -2500 -15687 2500 -15671
rect -2500 -15745 2500 -15729
rect -2500 -15779 -2484 -15745
rect 2484 -15779 2500 -15745
rect -2500 -15826 2500 -15779
rect -2500 -20873 2500 -20826
rect -2500 -20907 -2484 -20873
rect 2484 -20907 2500 -20873
rect -2500 -20923 2500 -20907
<< polycont >>
rect -2484 20873 2484 20907
rect -2484 15745 2484 15779
rect -2484 15637 2484 15671
rect -2484 10509 2484 10543
rect -2484 10401 2484 10435
rect -2484 5273 2484 5307
rect -2484 5165 2484 5199
rect -2484 37 2484 71
rect -2484 -71 2484 -37
rect -2484 -5199 2484 -5165
rect -2484 -5307 2484 -5273
rect -2484 -10435 2484 -10401
rect -2484 -10543 2484 -10509
rect -2484 -15671 2484 -15637
rect -2484 -15779 2484 -15745
rect -2484 -20907 2484 -20873
<< locali >>
rect -2660 20975 -2564 21009
rect 2564 20975 2660 21009
rect -2660 20913 -2626 20975
rect 2626 20913 2660 20975
rect -2500 20873 -2484 20907
rect 2484 20873 2500 20907
rect -2546 20814 -2512 20830
rect -2546 15822 -2512 15838
rect 2512 20814 2546 20830
rect 2512 15822 2546 15838
rect -2500 15745 -2484 15779
rect 2484 15745 2500 15779
rect -2500 15637 -2484 15671
rect 2484 15637 2500 15671
rect -2546 15578 -2512 15594
rect -2546 10586 -2512 10602
rect 2512 15578 2546 15594
rect 2512 10586 2546 10602
rect -2500 10509 -2484 10543
rect 2484 10509 2500 10543
rect -2500 10401 -2484 10435
rect 2484 10401 2500 10435
rect -2546 10342 -2512 10358
rect -2546 5350 -2512 5366
rect 2512 10342 2546 10358
rect 2512 5350 2546 5366
rect -2500 5273 -2484 5307
rect 2484 5273 2500 5307
rect -2500 5165 -2484 5199
rect 2484 5165 2500 5199
rect -2546 5106 -2512 5122
rect -2546 114 -2512 130
rect 2512 5106 2546 5122
rect 2512 114 2546 130
rect -2500 37 -2484 71
rect 2484 37 2500 71
rect -2500 -71 -2484 -37
rect 2484 -71 2500 -37
rect -2546 -130 -2512 -114
rect -2546 -5122 -2512 -5106
rect 2512 -130 2546 -114
rect 2512 -5122 2546 -5106
rect -2500 -5199 -2484 -5165
rect 2484 -5199 2500 -5165
rect -2500 -5307 -2484 -5273
rect 2484 -5307 2500 -5273
rect -2546 -5366 -2512 -5350
rect -2546 -10358 -2512 -10342
rect 2512 -5366 2546 -5350
rect 2512 -10358 2546 -10342
rect -2500 -10435 -2484 -10401
rect 2484 -10435 2500 -10401
rect -2500 -10543 -2484 -10509
rect 2484 -10543 2500 -10509
rect -2546 -10602 -2512 -10586
rect -2546 -15594 -2512 -15578
rect 2512 -10602 2546 -10586
rect 2512 -15594 2546 -15578
rect -2500 -15671 -2484 -15637
rect 2484 -15671 2500 -15637
rect -2500 -15779 -2484 -15745
rect 2484 -15779 2500 -15745
rect -2546 -15838 -2512 -15822
rect -2546 -20830 -2512 -20814
rect 2512 -15838 2546 -15822
rect 2512 -20830 2546 -20814
rect -2500 -20907 -2484 -20873
rect 2484 -20907 2500 -20873
rect -2660 -20975 -2626 -20913
rect 2626 -20975 2660 -20913
rect -2660 -21009 -2564 -20975
rect 2564 -21009 2660 -20975
<< viali >>
rect -2484 20873 2484 20907
rect -2546 15838 -2512 20814
rect 2512 15838 2546 20814
rect -2484 15745 2484 15779
rect -2484 15637 2484 15671
rect -2546 10602 -2512 15578
rect 2512 10602 2546 15578
rect -2484 10509 2484 10543
rect -2484 10401 2484 10435
rect -2546 5366 -2512 10342
rect 2512 5366 2546 10342
rect -2484 5273 2484 5307
rect -2484 5165 2484 5199
rect -2546 130 -2512 5106
rect 2512 130 2546 5106
rect -2484 37 2484 71
rect -2484 -71 2484 -37
rect -2546 -5106 -2512 -130
rect 2512 -5106 2546 -130
rect -2484 -5199 2484 -5165
rect -2484 -5307 2484 -5273
rect -2546 -10342 -2512 -5366
rect 2512 -10342 2546 -5366
rect -2484 -10435 2484 -10401
rect -2484 -10543 2484 -10509
rect -2546 -15578 -2512 -10602
rect 2512 -15578 2546 -10602
rect -2484 -15671 2484 -15637
rect -2484 -15779 2484 -15745
rect -2546 -20814 -2512 -15838
rect 2512 -20814 2546 -15838
rect -2484 -20907 2484 -20873
<< metal1 >>
rect -2496 20907 2496 20913
rect -2496 20873 -2484 20907
rect 2484 20873 2496 20907
rect -2496 20867 2496 20873
rect -2552 20814 -2506 20826
rect -2552 15838 -2546 20814
rect -2512 15838 -2506 20814
rect -2552 15826 -2506 15838
rect 2506 20814 2552 20826
rect 2506 15838 2512 20814
rect 2546 15838 2552 20814
rect 2506 15826 2552 15838
rect -2496 15779 2496 15785
rect -2496 15745 -2484 15779
rect 2484 15745 2496 15779
rect -2496 15739 2496 15745
rect -2496 15671 2496 15677
rect -2496 15637 -2484 15671
rect 2484 15637 2496 15671
rect -2496 15631 2496 15637
rect -2552 15578 -2506 15590
rect -2552 10602 -2546 15578
rect -2512 10602 -2506 15578
rect -2552 10590 -2506 10602
rect 2506 15578 2552 15590
rect 2506 10602 2512 15578
rect 2546 10602 2552 15578
rect 2506 10590 2552 10602
rect -2496 10543 2496 10549
rect -2496 10509 -2484 10543
rect 2484 10509 2496 10543
rect -2496 10503 2496 10509
rect -2496 10435 2496 10441
rect -2496 10401 -2484 10435
rect 2484 10401 2496 10435
rect -2496 10395 2496 10401
rect -2552 10342 -2506 10354
rect -2552 5366 -2546 10342
rect -2512 5366 -2506 10342
rect -2552 5354 -2506 5366
rect 2506 10342 2552 10354
rect 2506 5366 2512 10342
rect 2546 5366 2552 10342
rect 2506 5354 2552 5366
rect -2496 5307 2496 5313
rect -2496 5273 -2484 5307
rect 2484 5273 2496 5307
rect -2496 5267 2496 5273
rect -2496 5199 2496 5205
rect -2496 5165 -2484 5199
rect 2484 5165 2496 5199
rect -2496 5159 2496 5165
rect -2552 5106 -2506 5118
rect -2552 130 -2546 5106
rect -2512 130 -2506 5106
rect -2552 118 -2506 130
rect 2506 5106 2552 5118
rect 2506 130 2512 5106
rect 2546 130 2552 5106
rect 2506 118 2552 130
rect -2496 71 2496 77
rect -2496 37 -2484 71
rect 2484 37 2496 71
rect -2496 31 2496 37
rect -2496 -37 2496 -31
rect -2496 -71 -2484 -37
rect 2484 -71 2496 -37
rect -2496 -77 2496 -71
rect -2552 -130 -2506 -118
rect -2552 -5106 -2546 -130
rect -2512 -5106 -2506 -130
rect -2552 -5118 -2506 -5106
rect 2506 -130 2552 -118
rect 2506 -5106 2512 -130
rect 2546 -5106 2552 -130
rect 2506 -5118 2552 -5106
rect -2496 -5165 2496 -5159
rect -2496 -5199 -2484 -5165
rect 2484 -5199 2496 -5165
rect -2496 -5205 2496 -5199
rect -2496 -5273 2496 -5267
rect -2496 -5307 -2484 -5273
rect 2484 -5307 2496 -5273
rect -2496 -5313 2496 -5307
rect -2552 -5366 -2506 -5354
rect -2552 -10342 -2546 -5366
rect -2512 -10342 -2506 -5366
rect -2552 -10354 -2506 -10342
rect 2506 -5366 2552 -5354
rect 2506 -10342 2512 -5366
rect 2546 -10342 2552 -5366
rect 2506 -10354 2552 -10342
rect -2496 -10401 2496 -10395
rect -2496 -10435 -2484 -10401
rect 2484 -10435 2496 -10401
rect -2496 -10441 2496 -10435
rect -2496 -10509 2496 -10503
rect -2496 -10543 -2484 -10509
rect 2484 -10543 2496 -10509
rect -2496 -10549 2496 -10543
rect -2552 -10602 -2506 -10590
rect -2552 -15578 -2546 -10602
rect -2512 -15578 -2506 -10602
rect -2552 -15590 -2506 -15578
rect 2506 -10602 2552 -10590
rect 2506 -15578 2512 -10602
rect 2546 -15578 2552 -10602
rect 2506 -15590 2552 -15578
rect -2496 -15637 2496 -15631
rect -2496 -15671 -2484 -15637
rect 2484 -15671 2496 -15637
rect -2496 -15677 2496 -15671
rect -2496 -15745 2496 -15739
rect -2496 -15779 -2484 -15745
rect 2484 -15779 2496 -15745
rect -2496 -15785 2496 -15779
rect -2552 -15838 -2506 -15826
rect -2552 -20814 -2546 -15838
rect -2512 -20814 -2506 -15838
rect -2552 -20826 -2506 -20814
rect 2506 -15838 2552 -15826
rect 2506 -20814 2512 -15838
rect 2546 -20814 2552 -15838
rect 2506 -20826 2552 -20814
rect -2496 -20873 2496 -20867
rect -2496 -20907 -2484 -20873
rect 2484 -20907 2496 -20873
rect -2496 -20913 2496 -20907
<< labels >>
rlabel nsubdiffcont 0 -20992 0 -20992 0 B
port 1 nsew
rlabel pdiffc -2529 -18326 -2529 -18326 0 D0
port 2 nsew
rlabel pdiffc 2529 -18326 2529 -18326 0 S0
port 3 nsew
rlabel polycont 0 -15762 0 -15762 0 G0
port 4 nsew
rlabel pdiffc -2529 -13090 -2529 -13090 0 D1
port 5 nsew
rlabel pdiffc 2529 -13090 2529 -13090 0 S1
port 6 nsew
rlabel polycont 0 -10526 0 -10526 0 G1
port 7 nsew
rlabel pdiffc -2529 -7854 -2529 -7854 0 D2
port 8 nsew
rlabel pdiffc 2529 -7854 2529 -7854 0 S2
port 9 nsew
rlabel polycont 0 -5290 0 -5290 0 G2
port 10 nsew
rlabel pdiffc -2529 -2618 -2529 -2618 0 D3
port 11 nsew
rlabel pdiffc 2529 -2618 2529 -2618 0 S3
port 12 nsew
rlabel polycont 0 -54 0 -54 0 G3
port 13 nsew
rlabel pdiffc -2529 2618 -2529 2618 0 D4
port 14 nsew
rlabel pdiffc 2529 2618 2529 2618 0 S4
port 15 nsew
rlabel polycont 0 5182 0 5182 0 G4
port 16 nsew
rlabel pdiffc -2529 7854 -2529 7854 0 D5
port 17 nsew
rlabel pdiffc 2529 7854 2529 7854 0 S5
port 18 nsew
rlabel polycont 0 10418 0 10418 0 G5
port 19 nsew
rlabel pdiffc -2529 13090 -2529 13090 0 D6
port 20 nsew
rlabel pdiffc 2529 13090 2529 13090 0 S6
port 21 nsew
rlabel polycont 0 15654 0 15654 0 G6
port 22 nsew
rlabel pdiffc -2529 18326 -2529 18326 0 D7
port 23 nsew
rlabel pdiffc 2529 18326 2529 18326 0 S7
port 24 nsew
rlabel polycont 0 20890 0 20890 0 G7
port 25 nsew
<< properties >>
string FIXED_BBOX -2643 -20992 2643 20992
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 25.0 l 25.0 m 8 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
