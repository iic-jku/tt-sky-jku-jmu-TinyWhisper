magic
tech sky130A
magscale 1 2
timestamp 1762704370
<< metal3 >>
rect -3912 3312 -2880 3340
rect -3912 2688 -2964 3312
rect -2900 2688 -2880 3312
rect -3912 2660 -2880 2688
rect -2214 3312 -1182 3340
rect -2214 2688 -1266 3312
rect -1202 2688 -1182 3312
rect -2214 2660 -1182 2688
rect -516 3312 516 3340
rect -516 2688 432 3312
rect 496 2688 516 3312
rect -516 2660 516 2688
rect 1182 3312 2214 3340
rect 1182 2688 2130 3312
rect 2194 2688 2214 3312
rect 1182 2660 2214 2688
rect 2880 3312 3912 3340
rect 2880 2688 3828 3312
rect 3892 2688 3912 3312
rect 2880 2660 3912 2688
rect -3912 2312 -2880 2340
rect -3912 1688 -2964 2312
rect -2900 1688 -2880 2312
rect -3912 1660 -2880 1688
rect -2214 2312 -1182 2340
rect -2214 1688 -1266 2312
rect -1202 1688 -1182 2312
rect -2214 1660 -1182 1688
rect -516 2312 516 2340
rect -516 1688 432 2312
rect 496 1688 516 2312
rect -516 1660 516 1688
rect 1182 2312 2214 2340
rect 1182 1688 2130 2312
rect 2194 1688 2214 2312
rect 1182 1660 2214 1688
rect 2880 2312 3912 2340
rect 2880 1688 3828 2312
rect 3892 1688 3912 2312
rect 2880 1660 3912 1688
rect -3912 1312 -2880 1340
rect -3912 688 -2964 1312
rect -2900 688 -2880 1312
rect -3912 660 -2880 688
rect -2214 1312 -1182 1340
rect -2214 688 -1266 1312
rect -1202 688 -1182 1312
rect -2214 660 -1182 688
rect -516 1312 516 1340
rect -516 688 432 1312
rect 496 688 516 1312
rect -516 660 516 688
rect 1182 1312 2214 1340
rect 1182 688 2130 1312
rect 2194 688 2214 1312
rect 1182 660 2214 688
rect 2880 1312 3912 1340
rect 2880 688 3828 1312
rect 3892 688 3912 1312
rect 2880 660 3912 688
rect -3912 312 -2880 340
rect -3912 -312 -2964 312
rect -2900 -312 -2880 312
rect -3912 -340 -2880 -312
rect -2214 312 -1182 340
rect -2214 -312 -1266 312
rect -1202 -312 -1182 312
rect -2214 -340 -1182 -312
rect -516 312 516 340
rect -516 -312 432 312
rect 496 -312 516 312
rect -516 -340 516 -312
rect 1182 312 2214 340
rect 1182 -312 2130 312
rect 2194 -312 2214 312
rect 1182 -340 2214 -312
rect 2880 312 3912 340
rect 2880 -312 3828 312
rect 3892 -312 3912 312
rect 2880 -340 3912 -312
rect -3912 -688 -2880 -660
rect -3912 -1312 -2964 -688
rect -2900 -1312 -2880 -688
rect -3912 -1340 -2880 -1312
rect -2214 -688 -1182 -660
rect -2214 -1312 -1266 -688
rect -1202 -1312 -1182 -688
rect -2214 -1340 -1182 -1312
rect -516 -688 516 -660
rect -516 -1312 432 -688
rect 496 -1312 516 -688
rect -516 -1340 516 -1312
rect 1182 -688 2214 -660
rect 1182 -1312 2130 -688
rect 2194 -1312 2214 -688
rect 1182 -1340 2214 -1312
rect 2880 -688 3912 -660
rect 2880 -1312 3828 -688
rect 3892 -1312 3912 -688
rect 2880 -1340 3912 -1312
rect -3912 -1688 -2880 -1660
rect -3912 -2312 -2964 -1688
rect -2900 -2312 -2880 -1688
rect -3912 -2340 -2880 -2312
rect -2214 -1688 -1182 -1660
rect -2214 -2312 -1266 -1688
rect -1202 -2312 -1182 -1688
rect -2214 -2340 -1182 -2312
rect -516 -1688 516 -1660
rect -516 -2312 432 -1688
rect 496 -2312 516 -1688
rect -516 -2340 516 -2312
rect 1182 -1688 2214 -1660
rect 1182 -2312 2130 -1688
rect 2194 -2312 2214 -1688
rect 1182 -2340 2214 -2312
rect 2880 -1688 3912 -1660
rect 2880 -2312 3828 -1688
rect 3892 -2312 3912 -1688
rect 2880 -2340 3912 -2312
rect -3912 -2688 -2880 -2660
rect -3912 -3312 -2964 -2688
rect -2900 -3312 -2880 -2688
rect -3912 -3340 -2880 -3312
rect -2214 -2688 -1182 -2660
rect -2214 -3312 -1266 -2688
rect -1202 -3312 -1182 -2688
rect -2214 -3340 -1182 -3312
rect -516 -2688 516 -2660
rect -516 -3312 432 -2688
rect 496 -3312 516 -2688
rect -516 -3340 516 -3312
rect 1182 -2688 2214 -2660
rect 1182 -3312 2130 -2688
rect 2194 -3312 2214 -2688
rect 1182 -3340 2214 -3312
rect 2880 -2688 3912 -2660
rect 2880 -3312 3828 -2688
rect 3892 -3312 3912 -2688
rect 2880 -3340 3912 -3312
<< via3 >>
rect -2964 2688 -2900 3312
rect -1266 2688 -1202 3312
rect 432 2688 496 3312
rect 2130 2688 2194 3312
rect 3828 2688 3892 3312
rect -2964 1688 -2900 2312
rect -1266 1688 -1202 2312
rect 432 1688 496 2312
rect 2130 1688 2194 2312
rect 3828 1688 3892 2312
rect -2964 688 -2900 1312
rect -1266 688 -1202 1312
rect 432 688 496 1312
rect 2130 688 2194 1312
rect 3828 688 3892 1312
rect -2964 -312 -2900 312
rect -1266 -312 -1202 312
rect 432 -312 496 312
rect 2130 -312 2194 312
rect 3828 -312 3892 312
rect -2964 -1312 -2900 -688
rect -1266 -1312 -1202 -688
rect 432 -1312 496 -688
rect 2130 -1312 2194 -688
rect 3828 -1312 3892 -688
rect -2964 -2312 -2900 -1688
rect -1266 -2312 -1202 -1688
rect 432 -2312 496 -1688
rect 2130 -2312 2194 -1688
rect 3828 -2312 3892 -1688
rect -2964 -3312 -2900 -2688
rect -1266 -3312 -1202 -2688
rect 432 -3312 496 -2688
rect 2130 -3312 2194 -2688
rect 3828 -3312 3892 -2688
<< mimcap >>
rect -3872 3260 -3272 3300
rect -3872 2740 -3832 3260
rect -3312 2740 -3272 3260
rect -3872 2700 -3272 2740
rect -2174 3260 -1574 3300
rect -2174 2740 -2134 3260
rect -1614 2740 -1574 3260
rect -2174 2700 -1574 2740
rect -476 3260 124 3300
rect -476 2740 -436 3260
rect 84 2740 124 3260
rect -476 2700 124 2740
rect 1222 3260 1822 3300
rect 1222 2740 1262 3260
rect 1782 2740 1822 3260
rect 1222 2700 1822 2740
rect 2920 3260 3520 3300
rect 2920 2740 2960 3260
rect 3480 2740 3520 3260
rect 2920 2700 3520 2740
rect -3872 2260 -3272 2300
rect -3872 1740 -3832 2260
rect -3312 1740 -3272 2260
rect -3872 1700 -3272 1740
rect -2174 2260 -1574 2300
rect -2174 1740 -2134 2260
rect -1614 1740 -1574 2260
rect -2174 1700 -1574 1740
rect -476 2260 124 2300
rect -476 1740 -436 2260
rect 84 1740 124 2260
rect -476 1700 124 1740
rect 1222 2260 1822 2300
rect 1222 1740 1262 2260
rect 1782 1740 1822 2260
rect 1222 1700 1822 1740
rect 2920 2260 3520 2300
rect 2920 1740 2960 2260
rect 3480 1740 3520 2260
rect 2920 1700 3520 1740
rect -3872 1260 -3272 1300
rect -3872 740 -3832 1260
rect -3312 740 -3272 1260
rect -3872 700 -3272 740
rect -2174 1260 -1574 1300
rect -2174 740 -2134 1260
rect -1614 740 -1574 1260
rect -2174 700 -1574 740
rect -476 1260 124 1300
rect -476 740 -436 1260
rect 84 740 124 1260
rect -476 700 124 740
rect 1222 1260 1822 1300
rect 1222 740 1262 1260
rect 1782 740 1822 1260
rect 1222 700 1822 740
rect 2920 1260 3520 1300
rect 2920 740 2960 1260
rect 3480 740 3520 1260
rect 2920 700 3520 740
rect -3872 260 -3272 300
rect -3872 -260 -3832 260
rect -3312 -260 -3272 260
rect -3872 -300 -3272 -260
rect -2174 260 -1574 300
rect -2174 -260 -2134 260
rect -1614 -260 -1574 260
rect -2174 -300 -1574 -260
rect -476 260 124 300
rect -476 -260 -436 260
rect 84 -260 124 260
rect -476 -300 124 -260
rect 1222 260 1822 300
rect 1222 -260 1262 260
rect 1782 -260 1822 260
rect 1222 -300 1822 -260
rect 2920 260 3520 300
rect 2920 -260 2960 260
rect 3480 -260 3520 260
rect 2920 -300 3520 -260
rect -3872 -740 -3272 -700
rect -3872 -1260 -3832 -740
rect -3312 -1260 -3272 -740
rect -3872 -1300 -3272 -1260
rect -2174 -740 -1574 -700
rect -2174 -1260 -2134 -740
rect -1614 -1260 -1574 -740
rect -2174 -1300 -1574 -1260
rect -476 -740 124 -700
rect -476 -1260 -436 -740
rect 84 -1260 124 -740
rect -476 -1300 124 -1260
rect 1222 -740 1822 -700
rect 1222 -1260 1262 -740
rect 1782 -1260 1822 -740
rect 1222 -1300 1822 -1260
rect 2920 -740 3520 -700
rect 2920 -1260 2960 -740
rect 3480 -1260 3520 -740
rect 2920 -1300 3520 -1260
rect -3872 -1740 -3272 -1700
rect -3872 -2260 -3832 -1740
rect -3312 -2260 -3272 -1740
rect -3872 -2300 -3272 -2260
rect -2174 -1740 -1574 -1700
rect -2174 -2260 -2134 -1740
rect -1614 -2260 -1574 -1740
rect -2174 -2300 -1574 -2260
rect -476 -1740 124 -1700
rect -476 -2260 -436 -1740
rect 84 -2260 124 -1740
rect -476 -2300 124 -2260
rect 1222 -1740 1822 -1700
rect 1222 -2260 1262 -1740
rect 1782 -2260 1822 -1740
rect 1222 -2300 1822 -2260
rect 2920 -1740 3520 -1700
rect 2920 -2260 2960 -1740
rect 3480 -2260 3520 -1740
rect 2920 -2300 3520 -2260
rect -3872 -2740 -3272 -2700
rect -3872 -3260 -3832 -2740
rect -3312 -3260 -3272 -2740
rect -3872 -3300 -3272 -3260
rect -2174 -2740 -1574 -2700
rect -2174 -3260 -2134 -2740
rect -1614 -3260 -1574 -2740
rect -2174 -3300 -1574 -3260
rect -476 -2740 124 -2700
rect -476 -3260 -436 -2740
rect 84 -3260 124 -2740
rect -476 -3300 124 -3260
rect 1222 -2740 1822 -2700
rect 1222 -3260 1262 -2740
rect 1782 -3260 1822 -2740
rect 1222 -3300 1822 -3260
rect 2920 -2740 3520 -2700
rect 2920 -3260 2960 -2740
rect 3480 -3260 3520 -2740
rect 2920 -3300 3520 -3260
<< mimcapcontact >>
rect -3832 2740 -3312 3260
rect -2134 2740 -1614 3260
rect -436 2740 84 3260
rect 1262 2740 1782 3260
rect 2960 2740 3480 3260
rect -3832 1740 -3312 2260
rect -2134 1740 -1614 2260
rect -436 1740 84 2260
rect 1262 1740 1782 2260
rect 2960 1740 3480 2260
rect -3832 740 -3312 1260
rect -2134 740 -1614 1260
rect -436 740 84 1260
rect 1262 740 1782 1260
rect 2960 740 3480 1260
rect -3832 -260 -3312 260
rect -2134 -260 -1614 260
rect -436 -260 84 260
rect 1262 -260 1782 260
rect 2960 -260 3480 260
rect -3832 -1260 -3312 -740
rect -2134 -1260 -1614 -740
rect -436 -1260 84 -740
rect 1262 -1260 1782 -740
rect 2960 -1260 3480 -740
rect -3832 -2260 -3312 -1740
rect -2134 -2260 -1614 -1740
rect -436 -2260 84 -1740
rect 1262 -2260 1782 -1740
rect 2960 -2260 3480 -1740
rect -3832 -3260 -3312 -2740
rect -2134 -3260 -1614 -2740
rect -436 -3260 84 -2740
rect 1262 -3260 1782 -2740
rect 2960 -3260 3480 -2740
<< metal4 >>
rect -3624 3261 -3520 3500
rect -2984 3312 -2880 3500
rect -3833 3260 -3311 3261
rect -3833 2740 -3832 3260
rect -3312 2740 -3311 3260
rect -3833 2739 -3311 2740
rect -3624 2261 -3520 2739
rect -2984 2688 -2964 3312
rect -2900 2688 -2880 3312
rect -1926 3261 -1822 3500
rect -1286 3312 -1182 3500
rect -2135 3260 -1613 3261
rect -2135 2740 -2134 3260
rect -1614 2740 -1613 3260
rect -2135 2739 -1613 2740
rect -2984 2312 -2880 2688
rect -3833 2260 -3311 2261
rect -3833 1740 -3832 2260
rect -3312 1740 -3311 2260
rect -3833 1739 -3311 1740
rect -3624 1261 -3520 1739
rect -2984 1688 -2964 2312
rect -2900 1688 -2880 2312
rect -1926 2261 -1822 2739
rect -1286 2688 -1266 3312
rect -1202 2688 -1182 3312
rect -228 3261 -124 3500
rect 412 3312 516 3500
rect -437 3260 85 3261
rect -437 2740 -436 3260
rect 84 2740 85 3260
rect -437 2739 85 2740
rect -1286 2312 -1182 2688
rect -2135 2260 -1613 2261
rect -2135 1740 -2134 2260
rect -1614 1740 -1613 2260
rect -2135 1739 -1613 1740
rect -2984 1312 -2880 1688
rect -3833 1260 -3311 1261
rect -3833 740 -3832 1260
rect -3312 740 -3311 1260
rect -3833 739 -3311 740
rect -3624 261 -3520 739
rect -2984 688 -2964 1312
rect -2900 688 -2880 1312
rect -1926 1261 -1822 1739
rect -1286 1688 -1266 2312
rect -1202 1688 -1182 2312
rect -228 2261 -124 2739
rect 412 2688 432 3312
rect 496 2688 516 3312
rect 1470 3261 1574 3500
rect 2110 3312 2214 3500
rect 1261 3260 1783 3261
rect 1261 2740 1262 3260
rect 1782 2740 1783 3260
rect 1261 2739 1783 2740
rect 412 2312 516 2688
rect -437 2260 85 2261
rect -437 1740 -436 2260
rect 84 1740 85 2260
rect -437 1739 85 1740
rect -1286 1312 -1182 1688
rect -2135 1260 -1613 1261
rect -2135 740 -2134 1260
rect -1614 740 -1613 1260
rect -2135 739 -1613 740
rect -2984 312 -2880 688
rect -3833 260 -3311 261
rect -3833 -260 -3832 260
rect -3312 -260 -3311 260
rect -3833 -261 -3311 -260
rect -3624 -739 -3520 -261
rect -2984 -312 -2964 312
rect -2900 -312 -2880 312
rect -1926 261 -1822 739
rect -1286 688 -1266 1312
rect -1202 688 -1182 1312
rect -228 1261 -124 1739
rect 412 1688 432 2312
rect 496 1688 516 2312
rect 1470 2261 1574 2739
rect 2110 2688 2130 3312
rect 2194 2688 2214 3312
rect 3168 3261 3272 3500
rect 3808 3312 3912 3500
rect 2959 3260 3481 3261
rect 2959 2740 2960 3260
rect 3480 2740 3481 3260
rect 2959 2739 3481 2740
rect 2110 2312 2214 2688
rect 1261 2260 1783 2261
rect 1261 1740 1262 2260
rect 1782 1740 1783 2260
rect 1261 1739 1783 1740
rect 412 1312 516 1688
rect -437 1260 85 1261
rect -437 740 -436 1260
rect 84 740 85 1260
rect -437 739 85 740
rect -1286 312 -1182 688
rect -2135 260 -1613 261
rect -2135 -260 -2134 260
rect -1614 -260 -1613 260
rect -2135 -261 -1613 -260
rect -2984 -688 -2880 -312
rect -3833 -740 -3311 -739
rect -3833 -1260 -3832 -740
rect -3312 -1260 -3311 -740
rect -3833 -1261 -3311 -1260
rect -3624 -1739 -3520 -1261
rect -2984 -1312 -2964 -688
rect -2900 -1312 -2880 -688
rect -1926 -739 -1822 -261
rect -1286 -312 -1266 312
rect -1202 -312 -1182 312
rect -228 261 -124 739
rect 412 688 432 1312
rect 496 688 516 1312
rect 1470 1261 1574 1739
rect 2110 1688 2130 2312
rect 2194 1688 2214 2312
rect 3168 2261 3272 2739
rect 3808 2688 3828 3312
rect 3892 2688 3912 3312
rect 3808 2312 3912 2688
rect 2959 2260 3481 2261
rect 2959 1740 2960 2260
rect 3480 1740 3481 2260
rect 2959 1739 3481 1740
rect 2110 1312 2214 1688
rect 1261 1260 1783 1261
rect 1261 740 1262 1260
rect 1782 740 1783 1260
rect 1261 739 1783 740
rect 412 312 516 688
rect -437 260 85 261
rect -437 -260 -436 260
rect 84 -260 85 260
rect -437 -261 85 -260
rect -1286 -688 -1182 -312
rect -2135 -740 -1613 -739
rect -2135 -1260 -2134 -740
rect -1614 -1260 -1613 -740
rect -2135 -1261 -1613 -1260
rect -2984 -1688 -2880 -1312
rect -3833 -1740 -3311 -1739
rect -3833 -2260 -3832 -1740
rect -3312 -2260 -3311 -1740
rect -3833 -2261 -3311 -2260
rect -3624 -2739 -3520 -2261
rect -2984 -2312 -2964 -1688
rect -2900 -2312 -2880 -1688
rect -1926 -1739 -1822 -1261
rect -1286 -1312 -1266 -688
rect -1202 -1312 -1182 -688
rect -228 -739 -124 -261
rect 412 -312 432 312
rect 496 -312 516 312
rect 1470 261 1574 739
rect 2110 688 2130 1312
rect 2194 688 2214 1312
rect 3168 1261 3272 1739
rect 3808 1688 3828 2312
rect 3892 1688 3912 2312
rect 3808 1312 3912 1688
rect 2959 1260 3481 1261
rect 2959 740 2960 1260
rect 3480 740 3481 1260
rect 2959 739 3481 740
rect 2110 312 2214 688
rect 1261 260 1783 261
rect 1261 -260 1262 260
rect 1782 -260 1783 260
rect 1261 -261 1783 -260
rect 412 -688 516 -312
rect -437 -740 85 -739
rect -437 -1260 -436 -740
rect 84 -1260 85 -740
rect -437 -1261 85 -1260
rect -1286 -1688 -1182 -1312
rect -2135 -1740 -1613 -1739
rect -2135 -2260 -2134 -1740
rect -1614 -2260 -1613 -1740
rect -2135 -2261 -1613 -2260
rect -2984 -2688 -2880 -2312
rect -3833 -2740 -3311 -2739
rect -3833 -3260 -3832 -2740
rect -3312 -3260 -3311 -2740
rect -3833 -3261 -3311 -3260
rect -3624 -3500 -3520 -3261
rect -2984 -3312 -2964 -2688
rect -2900 -3312 -2880 -2688
rect -1926 -2739 -1822 -2261
rect -1286 -2312 -1266 -1688
rect -1202 -2312 -1182 -1688
rect -228 -1739 -124 -1261
rect 412 -1312 432 -688
rect 496 -1312 516 -688
rect 1470 -739 1574 -261
rect 2110 -312 2130 312
rect 2194 -312 2214 312
rect 3168 261 3272 739
rect 3808 688 3828 1312
rect 3892 688 3912 1312
rect 3808 312 3912 688
rect 2959 260 3481 261
rect 2959 -260 2960 260
rect 3480 -260 3481 260
rect 2959 -261 3481 -260
rect 2110 -688 2214 -312
rect 1261 -740 1783 -739
rect 1261 -1260 1262 -740
rect 1782 -1260 1783 -740
rect 1261 -1261 1783 -1260
rect 412 -1688 516 -1312
rect -437 -1740 85 -1739
rect -437 -2260 -436 -1740
rect 84 -2260 85 -1740
rect -437 -2261 85 -2260
rect -1286 -2688 -1182 -2312
rect -2135 -2740 -1613 -2739
rect -2135 -3260 -2134 -2740
rect -1614 -3260 -1613 -2740
rect -2135 -3261 -1613 -3260
rect -2984 -3500 -2880 -3312
rect -1926 -3500 -1822 -3261
rect -1286 -3312 -1266 -2688
rect -1202 -3312 -1182 -2688
rect -228 -2739 -124 -2261
rect 412 -2312 432 -1688
rect 496 -2312 516 -1688
rect 1470 -1739 1574 -1261
rect 2110 -1312 2130 -688
rect 2194 -1312 2214 -688
rect 3168 -739 3272 -261
rect 3808 -312 3828 312
rect 3892 -312 3912 312
rect 3808 -688 3912 -312
rect 2959 -740 3481 -739
rect 2959 -1260 2960 -740
rect 3480 -1260 3481 -740
rect 2959 -1261 3481 -1260
rect 2110 -1688 2214 -1312
rect 1261 -1740 1783 -1739
rect 1261 -2260 1262 -1740
rect 1782 -2260 1783 -1740
rect 1261 -2261 1783 -2260
rect 412 -2688 516 -2312
rect -437 -2740 85 -2739
rect -437 -3260 -436 -2740
rect 84 -3260 85 -2740
rect -437 -3261 85 -3260
rect -1286 -3500 -1182 -3312
rect -228 -3500 -124 -3261
rect 412 -3312 432 -2688
rect 496 -3312 516 -2688
rect 1470 -2739 1574 -2261
rect 2110 -2312 2130 -1688
rect 2194 -2312 2214 -1688
rect 3168 -1739 3272 -1261
rect 3808 -1312 3828 -688
rect 3892 -1312 3912 -688
rect 3808 -1688 3912 -1312
rect 2959 -1740 3481 -1739
rect 2959 -2260 2960 -1740
rect 3480 -2260 3481 -1740
rect 2959 -2261 3481 -2260
rect 2110 -2688 2214 -2312
rect 1261 -2740 1783 -2739
rect 1261 -3260 1262 -2740
rect 1782 -3260 1783 -2740
rect 1261 -3261 1783 -3260
rect 412 -3500 516 -3312
rect 1470 -3500 1574 -3261
rect 2110 -3312 2130 -2688
rect 2194 -3312 2214 -2688
rect 3168 -2739 3272 -2261
rect 3808 -2312 3828 -1688
rect 3892 -2312 3912 -1688
rect 3808 -2688 3912 -2312
rect 2959 -2740 3481 -2739
rect 2959 -3260 2960 -2740
rect 3480 -3260 3481 -2740
rect 2959 -3261 3481 -3260
rect 2110 -3500 2214 -3312
rect 3168 -3500 3272 -3261
rect 3808 -3312 3828 -2688
rect 3892 -3312 3912 -2688
rect 3808 -3500 3912 -3312
<< labels >>
rlabel via3 -2932 -3000 -2932 -3000 0 C2_0
port 1 nsew
rlabel mimcapcontact -3572 -3000 -3572 -3000 0 C1_0
port 2 nsew
rlabel via3 -1234 -3000 -1234 -3000 0 C2_1
port 3 nsew
rlabel mimcapcontact -1874 -3000 -1874 -3000 0 C1_1
port 4 nsew
rlabel via3 464 -3000 464 -3000 0 C2_2
port 5 nsew
rlabel mimcapcontact -176 -3000 -176 -3000 0 C1_2
port 6 nsew
rlabel via3 2162 -3000 2162 -3000 0 C2_3
port 7 nsew
rlabel mimcapcontact 1522 -3000 1522 -3000 0 C1_3
port 8 nsew
rlabel via3 3860 -3000 3860 -3000 0 C2_4
port 9 nsew
rlabel mimcapcontact 3220 -3000 3220 -3000 0 C1_4
port 10 nsew
<< properties >>
string FIXED_BBOX 2880 2660 3560 3340
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 3.00 l 3.00 val 20.28 carea 2.00 cperi 0.19 class capacitor nx 5 ny 7 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100 stack 1 doports 1
<< end >>
