magic
tech sky130A
magscale 1 2
timestamp 1762641840
<< locali >>
rect 10 160 230 770
rect 760 160 980 770
rect 5 -520 230 -310
rect 760 -520 985 -310
<< viali >>
rect -40 180 0 750
rect 990 180 1030 750
rect -40 -500 0 -330
rect 990 -500 1030 -330
<< metal1 >>
rect -55 915 1045 985
rect -55 765 145 915
rect -55 750 190 765
rect -55 180 -40 750
rect 0 565 190 750
rect 270 755 335 765
rect 0 365 200 565
rect 0 180 190 365
rect -55 165 190 180
rect 270 175 275 755
rect 270 165 335 175
rect 375 165 425 915
rect 465 755 530 765
rect 465 175 470 755
rect 525 175 530 755
rect 465 165 530 175
rect 565 165 615 915
rect 845 765 1045 915
rect 655 755 720 765
rect 655 175 660 755
rect 715 175 720 755
rect 800 750 1045 765
rect 800 565 990 750
rect 795 365 990 565
rect 655 165 720 175
rect 800 180 990 365
rect 1030 180 1045 750
rect 800 165 1045 180
rect 220 -20 770 125
rect -70 -140 770 -20
rect 220 -275 770 -140
rect -55 -330 230 -315
rect -55 -500 -40 -330
rect 0 -500 230 -330
rect -55 -515 230 -500
rect 270 -325 335 -315
rect 270 -505 275 -325
rect 270 -515 335 -505
rect -55 -520 231 -515
rect -55 -655 230 -520
rect 375 -655 425 -315
rect 465 -325 530 -315
rect 465 -505 470 -325
rect 525 -505 530 -325
rect 465 -515 530 -505
rect 565 -655 615 -315
rect 655 -325 720 -315
rect 655 -505 660 -325
rect 715 -505 720 -325
rect 655 -515 720 -505
rect 760 -330 1045 -315
rect 760 -500 990 -330
rect 1030 -500 1045 -330
rect 760 -655 1045 -500
rect -55 -700 1045 -655
rect -55 -725 230 -700
rect 420 -720 570 -700
rect 760 -725 1045 -700
<< via1 >>
rect 275 175 335 755
rect 470 175 525 755
rect 660 175 715 755
rect 275 -505 335 -325
rect 470 -505 525 -325
rect 660 -505 715 -325
<< metal2 >>
rect 270 755 335 765
rect 270 175 275 755
rect 270 -20 335 175
rect 465 755 530 765
rect 465 175 470 755
rect 525 175 530 755
rect 465 -20 530 175
rect 655 755 720 765
rect 655 175 660 755
rect 715 175 720 755
rect 655 -20 720 175
rect 270 -140 1060 -20
rect 270 -325 335 -140
rect 270 -505 275 -325
rect 270 -515 335 -505
rect 465 -325 530 -140
rect 465 -505 470 -325
rect 525 -505 530 -325
rect 465 -515 530 -505
rect 655 -325 720 -140
rect 655 -505 660 -325
rect 715 -505 720 -325
rect 655 -515 720 -505
use sky130_fd_pr__nfet_01v8_4FXFJ2  sky130_fd_pr__nfet_01v8_4FXFJ2_0
timestamp 1762641840
transform 1 0 496 0 1 -415
box -551 -310 551 310
use sky130_fd_pr__pfet_01v8_JBT5N5  sky130_fd_pr__pfet_01v8_JBT5N5_0
timestamp 1762641840
transform 1 0 496 0 1 465
box -551 -520 551 520
<< labels >>
flabel metal1 -60 -80 -60 -80 0 FreeSans 400 0 0 0 vin
port 5 nsew
flabel metal1 495 950 495 950 0 FreeSans 400 0 0 0 VDD
port 13 nsew
flabel metal2 1050 -85 1050 -85 0 FreeSans 400 0 0 0 vout
port 15 nsew
flabel metal1 495 -690 495 -690 0 FreeSans 400 0 0 0 VSS
port 17 nsew
<< end >>
