magic
tech sky130A
magscale 1 2
timestamp 1762641840
<< nwell >>
rect -551 -519 551 519
<< pmos >>
rect -351 -300 -321 300
rect -255 -300 -225 300
rect -159 -300 -129 300
rect -63 -300 -33 300
rect 33 -300 63 300
rect 129 -300 159 300
rect 225 -300 255 300
rect 321 -300 351 300
<< pdiff >>
rect -413 288 -351 300
rect -413 -288 -401 288
rect -367 -288 -351 288
rect -413 -300 -351 -288
rect -321 288 -255 300
rect -321 -288 -305 288
rect -271 -288 -255 288
rect -321 -300 -255 -288
rect -225 288 -159 300
rect -225 -288 -209 288
rect -175 -288 -159 288
rect -225 -300 -159 -288
rect -129 288 -63 300
rect -129 -288 -113 288
rect -79 -288 -63 288
rect -129 -300 -63 -288
rect -33 288 33 300
rect -33 -288 -17 288
rect 17 -288 33 288
rect -33 -300 33 -288
rect 63 288 129 300
rect 63 -288 79 288
rect 113 -288 129 288
rect 63 -300 129 -288
rect 159 288 225 300
rect 159 -288 175 288
rect 209 -288 225 288
rect 159 -300 225 -288
rect 255 288 321 300
rect 255 -288 271 288
rect 305 -288 321 288
rect 255 -300 321 -288
rect 351 288 413 300
rect 351 -288 367 288
rect 401 -288 413 288
rect 351 -300 413 -288
<< pdiffc >>
rect -401 -288 -367 288
rect -305 -288 -271 288
rect -209 -288 -175 288
rect -113 -288 -79 288
rect -17 -288 17 288
rect 79 -288 113 288
rect 175 -288 209 288
rect 271 -288 305 288
rect 367 -288 401 288
<< nsubdiff >>
rect -515 449 -419 483
rect 419 449 515 483
rect -515 387 -481 449
rect 481 387 515 449
rect -515 -449 -481 -387
rect 481 -449 515 -387
rect -515 -483 -419 -449
rect 419 -483 515 -449
<< nsubdiffcont >>
rect -419 449 419 483
rect -515 -387 -481 387
rect 481 -387 515 387
rect -419 -483 419 -449
<< poly >>
rect -425 395 -321 415
rect -425 360 -405 395
rect -345 360 -321 395
rect -425 340 -321 360
rect -351 300 -321 340
rect 321 395 425 415
rect 321 360 345 395
rect 405 360 425 395
rect 321 340 425 360
rect -255 300 -225 326
rect -159 300 -129 326
rect -63 300 -33 326
rect 33 300 63 326
rect 129 300 159 326
rect 225 300 255 326
rect 321 300 351 340
rect -351 -326 -321 -300
rect -255 -340 -225 -300
rect -159 -340 -129 -300
rect -63 -340 -33 -300
rect 33 -340 63 -300
rect 129 -340 159 -300
rect 225 -340 255 -300
rect 321 -326 351 -300
rect -275 -360 275 -340
rect -275 -395 -255 -360
rect 255 -395 275 -360
rect -275 -415 275 -395
<< polycont >>
rect -405 360 -345 395
rect 345 360 405 395
rect -255 -395 255 -360
<< locali >>
rect -550 505 550 520
rect -550 465 -535 505
rect 535 465 550 505
rect -550 449 -419 465
rect 419 449 550 465
rect -550 387 -480 449
rect -550 -387 -515 387
rect -481 -387 -480 387
rect -425 400 -325 410
rect -425 355 -410 400
rect -365 395 -325 400
rect -345 360 -325 395
rect -365 355 -325 360
rect -425 345 -325 355
rect 325 400 425 410
rect 325 395 365 400
rect 325 360 345 395
rect 325 355 365 360
rect 410 355 425 400
rect 325 345 425 355
rect 480 387 550 449
rect -401 288 -367 304
rect -401 -304 -367 -288
rect -305 288 -271 304
rect -305 -304 -271 -288
rect -209 288 -175 304
rect -209 -304 -175 -288
rect -113 288 -79 304
rect -113 -304 -79 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 79 288 113 304
rect 79 -304 113 -288
rect 175 288 209 304
rect 175 -304 209 -288
rect 271 288 305 304
rect 271 -304 305 -288
rect 367 288 401 304
rect 367 -304 401 -288
rect -550 -449 -480 -387
rect -275 -355 275 -340
rect -275 -400 -260 -355
rect 260 -400 275 -355
rect -275 -415 275 -400
rect 480 -387 481 387
rect 515 -387 550 387
rect 480 -449 550 -387
rect -550 -483 -419 -449
rect 419 -483 550 -449
rect -550 -520 550 -483
<< viali >>
rect -535 483 535 505
rect -535 465 -419 483
rect -419 465 419 483
rect 419 465 535 483
rect -410 395 -365 400
rect -410 360 -405 395
rect -405 360 -365 395
rect -410 355 -365 360
rect 365 395 410 400
rect 365 360 405 395
rect 405 360 410 395
rect 365 355 410 360
rect -401 -288 -367 288
rect -305 -288 -271 288
rect -209 -288 -175 288
rect -113 -288 -79 288
rect -17 -288 17 288
rect 79 -288 113 288
rect 175 -288 209 288
rect 271 -288 305 288
rect 367 -288 401 288
rect -260 -360 260 -355
rect -260 -395 -255 -360
rect -255 -395 255 -360
rect 255 -395 260 -360
rect -260 -400 260 -395
<< metal1 >>
rect -550 505 550 520
rect -550 465 -535 505
rect 535 465 550 505
rect -550 450 550 465
rect -425 400 -350 410
rect -425 355 -410 400
rect -365 355 -350 400
rect -425 345 -350 355
rect 350 400 425 410
rect 350 355 365 400
rect 410 355 425 400
rect 350 345 425 355
rect -407 288 -361 300
rect -407 -288 -401 288
rect -367 -288 -361 288
rect -407 -300 -361 -288
rect -311 288 -265 300
rect -311 -288 -305 288
rect -271 -288 -265 288
rect -311 -300 -265 -288
rect -215 288 -169 300
rect -215 -288 -209 288
rect -175 -288 -169 288
rect -215 -300 -169 -288
rect -119 288 -73 300
rect -119 -288 -113 288
rect -79 -288 -73 288
rect -119 -300 -73 -288
rect -23 288 23 300
rect -23 -288 -17 288
rect 17 -288 23 288
rect -23 -300 23 -288
rect 73 288 119 300
rect 73 -288 79 288
rect 113 -288 119 288
rect 73 -300 119 -288
rect 169 288 215 300
rect 169 -288 175 288
rect 209 -288 215 288
rect 169 -300 215 -288
rect 265 288 311 300
rect 265 -288 271 288
rect 305 -288 311 288
rect 265 -300 311 -288
rect 361 288 407 300
rect 361 -288 367 288
rect 401 -288 407 288
rect 361 -300 407 -288
rect -275 -355 275 -340
rect -275 -400 -260 -355
rect 260 -400 275 -355
rect -275 -415 275 -400
<< labels >>
rlabel nsubdiffcont 0 -466 0 -466 0 B
port 1 nsew
rlabel pdiffc -384 0 -384 0 0 D0
port 2 nsew
rlabel pdiffc -288 0 -288 0 0 S1
port 4 nsew
rlabel pdiffc -192 0 -192 0 0 D2
port 6 nsew
rlabel pdiffc -96 0 -96 0 0 S3
port 8 nsew
rlabel pdiffc 0 0 0 0 0 D4
port 10 nsew
rlabel pdiffc 96 0 96 0 0 S5
port 12 nsew
rlabel pdiffc 192 0 192 0 0 D6
port 14 nsew
rlabel pdiffc 288 0 288 0 0 S7
port 16 nsew
<< properties >>
string FIXED_BBOX -498 -466 498 466
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3.0 l 0.15 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
