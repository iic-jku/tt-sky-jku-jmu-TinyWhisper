magic
tech sky130A
magscale 1 2
timestamp 1757014995
<< viali >>
rect -100 2290 -60 4065
rect 1680 2290 1720 4065
rect -100 1220 -60 1800
rect 1680 1220 1720 1800
<< metal1 >>
rect -130 4545 1755 4695
rect -130 4085 -25 4545
rect 70 4435 240 4450
rect 70 4315 85 4435
rect 225 4315 240 4435
rect 70 4130 240 4315
rect 1370 4435 1540 4450
rect 1370 4315 1385 4435
rect 1525 4315 1540 4435
rect 290 4135 1330 4170
rect -130 4065 240 4085
rect -130 2290 -100 4065
rect -60 2290 85 4065
rect 225 2290 240 4065
rect -130 2275 240 2290
rect 290 2275 325 4135
rect 500 4065 605 4080
rect 500 2290 515 4065
rect 590 2290 605 4065
rect 500 2275 605 2290
rect 795 2280 830 4135
rect 1015 4065 1120 4080
rect 1015 2290 1030 4065
rect 1105 2290 1120 4065
rect 1015 2275 1120 2290
rect 1295 2280 1330 4135
rect 1370 4130 1540 4315
rect 1650 4085 1755 4545
rect 1570 4065 1755 4085
rect 1570 2290 1680 4065
rect 1720 2290 1755 4065
rect 1570 2275 1755 2290
rect 330 2095 1300 2230
rect -165 1985 1300 2095
rect 330 1850 1300 1985
rect -130 1800 55 1815
rect -130 1220 -100 1800
rect -60 1220 55 1800
rect -130 1205 55 1220
rect -130 755 -25 1205
rect 70 985 240 1170
rect 290 1155 325 1810
rect 505 1795 595 1810
rect 505 1225 520 1795
rect 580 1225 595 1795
rect 505 1210 595 1225
rect 795 1155 830 1810
rect 1025 1795 1115 1810
rect 1025 1225 1040 1795
rect 1100 1225 1115 1795
rect 1025 1210 1115 1225
rect 1295 1155 1330 1810
rect 1570 1800 1755 1815
rect 1570 1220 1680 1800
rect 1720 1220 1755 1800
rect 1570 1205 1755 1220
rect 290 1120 1330 1155
rect 70 865 85 985
rect 225 865 240 985
rect 70 850 240 865
rect 1370 985 1540 1170
rect 1370 865 1385 985
rect 1525 865 1540 985
rect 1370 850 1540 865
rect 1650 755 1755 1205
rect -130 605 1755 755
<< via1 >>
rect 85 4315 225 4435
rect 1385 4315 1525 4435
rect 85 2290 225 4065
rect 515 2290 590 4065
rect 1030 2290 1105 4065
rect 520 1225 580 1795
rect 1040 1225 1100 1795
rect 85 865 225 985
rect 1385 865 1525 985
<< metal2 >>
rect -165 4435 1540 4450
rect -165 4315 85 4435
rect 225 4315 1385 4435
rect 1525 4315 1540 4435
rect -165 4300 1540 4315
rect 70 4065 240 4085
rect 70 2290 85 4065
rect 225 2290 240 4065
rect 70 1000 240 2290
rect 500 4065 605 4080
rect 500 2290 515 4065
rect 590 2290 605 4065
rect 500 2275 605 2290
rect 1015 4065 1120 4080
rect 1015 2290 1030 4065
rect 1105 2290 1120 4065
rect 1015 2275 1120 2290
rect 530 2095 575 2275
rect 1045 2095 1090 2275
rect 530 1985 1770 2095
rect 530 1810 575 1985
rect 1045 1810 1090 1985
rect 505 1795 595 1810
rect 505 1225 520 1795
rect 580 1225 595 1795
rect 505 1210 595 1225
rect 1025 1795 1115 1810
rect 1025 1225 1040 1795
rect 1100 1225 1115 1795
rect 1025 1210 1115 1225
rect 70 985 1540 1000
rect 70 865 85 985
rect 225 865 1385 985
rect 1525 865 1540 985
rect 70 850 1540 865
use sky130_fd_pr__nfet_01v8_lvt_XCBGUP  sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0
timestamp 1757014995
transform 1 0 811 0 1 1510
box -941 -510 941 510
use sky130_fd_pr__pfet_01v8_lvt_P4JB26  sky130_fd_pr__pfet_01v8_lvt_P4JB26_0
timestamp 1757014995
transform 1 0 811 0 1 3179
box -941 -1119 941 1119
<< labels >>
flabel metal2 -155 4370 -155 4370 0 FreeSans 320 0 0 0 di_en
port 8 nsew
flabel metal1 1040 670 1040 670 0 FreeSans 400 0 0 0 VSS
port 10 nsew
flabel metal1 965 4610 965 4610 0 FreeSans 400 0 0 0 VDD
port 11 nsew
flabel metal1 -155 2040 -155 2040 0 FreeSans 320 0 0 0 vin
port 12 nsew
flabel metal2 1760 2040 1760 2040 0 FreeSans 320 0 0 0 vout
port 14 nsew
<< end >>
