magic
tech sky130A
magscale 1 2
timestamp 1762641840
<< locali >>
rect -15 975 2910 990
rect -15 935 0 975
rect 2895 935 2910 975
rect -15 20 55 935
rect 2840 20 2910 935
rect -15 -50 2910 20
rect -15 -170 2910 -100
rect -15 -650 55 -170
rect 2840 -650 2910 -170
rect -15 -665 2910 -650
rect -15 -705 0 -665
rect 2895 -705 2910 -665
rect -15 -720 2910 -705
<< viali >>
rect 0 935 2895 975
rect 0 -705 2895 -665
<< metal1 >>
rect -15 975 2910 990
rect -15 935 0 975
rect 2895 935 2910 975
rect -15 920 2910 935
rect -15 810 2910 885
rect -15 -550 55 810
rect 120 745 560 755
rect 120 530 130 745
rect 460 530 560 745
rect 120 520 560 530
rect 600 745 665 755
rect 600 530 605 745
rect 660 530 665 745
rect 600 520 665 530
rect 790 745 855 755
rect 790 530 795 745
rect 850 530 855 745
rect 790 520 855 530
rect 985 745 1050 755
rect 985 530 990 745
rect 1045 530 1050 745
rect 985 520 1050 530
rect 1175 745 1240 755
rect 1175 530 1180 745
rect 1235 530 1240 745
rect 1175 520 1240 530
rect 1365 745 1435 755
rect 1365 530 1370 745
rect 1430 530 1435 745
rect 1365 520 1435 530
rect 1560 745 1625 755
rect 1560 530 1565 745
rect 1620 530 1625 745
rect 1560 520 1625 530
rect 1750 745 1815 755
rect 1750 530 1755 745
rect 1810 530 1815 745
rect 1750 520 1815 530
rect 1945 745 2010 755
rect 1945 530 1950 745
rect 2005 530 2010 745
rect 1945 520 2010 530
rect 2135 745 2200 755
rect 2135 530 2140 745
rect 2195 530 2200 745
rect 2135 520 2200 530
rect 2325 745 2775 755
rect 2325 530 2335 745
rect 2765 530 2775 745
rect 2325 520 2775 530
rect 505 405 515 520
rect 555 515 560 520
rect 555 405 570 515
rect 505 395 570 405
rect 505 180 510 395
rect 565 180 570 395
rect 505 170 570 180
rect 695 395 760 405
rect 695 180 700 395
rect 755 180 760 395
rect 695 170 760 180
rect 885 395 955 405
rect 885 180 890 395
rect 950 180 955 395
rect 885 170 955 180
rect 1080 395 1145 405
rect 1080 180 1085 395
rect 1140 180 1145 395
rect 1080 170 1145 180
rect 1270 395 1335 405
rect 1270 180 1275 395
rect 1330 180 1335 395
rect 1270 170 1335 180
rect 1465 395 1530 405
rect 1465 180 1470 395
rect 1525 180 1530 395
rect 1465 170 1530 180
rect 1655 395 1720 405
rect 1655 180 1660 395
rect 1715 180 1720 395
rect 1655 170 1720 180
rect 1845 395 1910 405
rect 1845 180 1850 395
rect 1905 180 1910 395
rect 1845 170 1910 180
rect 2040 395 2105 405
rect 2040 180 2045 395
rect 2100 180 2105 395
rect 2040 170 2105 180
rect 2230 395 2295 405
rect 2230 180 2235 395
rect 2230 170 2295 180
rect 165 -270 2730 130
rect 505 -320 570 -310
rect 505 -380 510 -320
rect 565 -380 570 -320
rect 505 -435 570 -380
rect 695 -320 760 -310
rect 695 -380 700 -320
rect 755 -380 760 -320
rect 695 -390 760 -380
rect 885 -320 955 -310
rect 885 -380 890 -320
rect 950 -380 955 -320
rect 885 -390 955 -380
rect 1080 -320 1145 -310
rect 1080 -380 1085 -320
rect 1140 -380 1145 -320
rect 1080 -390 1145 -380
rect 1270 -320 1335 -310
rect 1270 -380 1275 -320
rect 1330 -380 1335 -320
rect 1270 -390 1335 -380
rect 1465 -320 1530 -310
rect 1465 -380 1470 -320
rect 1525 -380 1530 -320
rect 1465 -390 1530 -380
rect 1655 -320 1720 -310
rect 1655 -380 1660 -320
rect 1715 -380 1720 -320
rect 1655 -390 1720 -380
rect 1845 -320 1915 -310
rect 1845 -380 1850 -320
rect 1910 -380 1915 -320
rect 1845 -390 1915 -380
rect 2040 -320 2105 -310
rect 2040 -380 2045 -320
rect 2100 -380 2105 -320
rect 2040 -390 2105 -380
rect 2230 -320 2300 -310
rect 2230 -380 2235 -320
rect 2295 -380 2300 -320
rect 2230 -390 2300 -380
rect 505 -440 565 -435
rect 120 -450 565 -440
rect 120 -510 130 -450
rect 460 -510 565 -450
rect 120 -520 565 -510
rect 600 -450 665 -440
rect 600 -510 605 -450
rect 660 -510 665 -450
rect 600 -520 665 -510
rect 790 -450 860 -440
rect 790 -510 795 -450
rect 850 -510 860 -450
rect 790 -520 860 -510
rect 985 -450 1050 -440
rect 985 -510 990 -450
rect 1045 -510 1050 -450
rect 985 -520 1050 -510
rect 1175 -450 1240 -440
rect 1175 -510 1180 -450
rect 1235 -510 1240 -450
rect 1175 -520 1240 -510
rect 1365 -450 1435 -440
rect 1365 -510 1375 -450
rect 1430 -510 1435 -450
rect 1365 -520 1435 -510
rect 1560 -450 1625 -440
rect 1560 -510 1565 -450
rect 1620 -510 1625 -450
rect 1560 -520 1625 -510
rect 1750 -450 1820 -440
rect 1750 -510 1755 -450
rect 1810 -510 1820 -450
rect 1750 -520 1820 -510
rect 1945 -450 2010 -440
rect 1945 -510 1950 -450
rect 2005 -510 2010 -450
rect 1945 -520 2010 -510
rect 2135 -450 2200 -440
rect 2135 -510 2140 -450
rect 2195 -510 2200 -450
rect 2135 -520 2200 -510
rect 2325 -450 2775 -440
rect 2325 -510 2340 -450
rect 2765 -510 2775 -450
rect 2325 -520 2775 -510
rect 2840 -550 2910 810
rect -15 -615 560 -550
rect 2340 -615 2910 -550
rect -15 -665 2910 -650
rect -15 -705 0 -665
rect 2895 -705 2910 -665
rect -15 -720 2910 -705
<< via1 >>
rect 130 530 460 745
rect 605 530 660 745
rect 795 530 850 745
rect 990 530 1045 745
rect 1180 530 1235 745
rect 1370 530 1430 745
rect 1565 530 1620 745
rect 1755 530 1810 745
rect 1950 530 2005 745
rect 2140 530 2195 745
rect 2335 530 2765 745
rect 510 180 565 395
rect 700 180 755 395
rect 890 180 950 395
rect 1085 180 1140 395
rect 1275 180 1330 395
rect 1470 180 1525 395
rect 1660 180 1715 395
rect 1850 180 1905 395
rect 2045 180 2100 395
rect 2235 180 2295 395
rect 510 -380 565 -320
rect 700 -380 755 -320
rect 890 -380 950 -320
rect 1085 -380 1140 -320
rect 1275 -380 1330 -320
rect 1470 -380 1525 -320
rect 1660 -380 1715 -320
rect 1850 -380 1910 -320
rect 2045 -380 2100 -320
rect 2235 -380 2295 -320
rect 130 -510 460 -450
rect 605 -510 660 -450
rect 795 -510 850 -450
rect 990 -510 1045 -450
rect 1180 -510 1235 -450
rect 1375 -510 1430 -450
rect 1565 -510 1620 -450
rect 1755 -510 1810 -450
rect 1950 -510 2005 -450
rect 2140 -510 2195 -450
rect 2340 -510 2765 -450
<< metal2 >>
rect 120 745 470 755
rect 120 530 130 745
rect 460 530 470 745
rect 120 520 470 530
rect 600 745 2775 755
rect 600 530 605 745
rect 660 530 795 745
rect 850 530 990 745
rect 1045 530 1180 745
rect 1235 530 1370 745
rect 1430 530 1565 745
rect 1620 530 1755 745
rect 1810 530 1950 745
rect 2005 530 2140 745
rect 2195 530 2335 745
rect 2765 530 2775 745
rect 600 520 2775 530
rect 500 180 510 395
rect 565 180 700 395
rect 755 180 890 395
rect 950 180 1085 395
rect 1140 180 1275 395
rect 1330 180 1470 395
rect 1525 180 1660 395
rect 1715 180 1850 395
rect 1905 180 2045 395
rect 2100 180 2235 395
rect 2295 180 2305 395
rect 500 -320 2305 180
rect 500 -380 510 -320
rect 565 -380 700 -320
rect 755 -380 890 -320
rect 950 -380 1085 -320
rect 1140 -380 1275 -320
rect 1330 -380 1470 -320
rect 1525 -380 1660 -320
rect 1715 -380 1850 -320
rect 1910 -380 2045 -320
rect 2100 -380 2235 -320
rect 2295 -380 2305 -320
rect 120 -450 465 -440
rect 120 -510 130 -450
rect 460 -510 465 -450
rect 120 -520 465 -510
rect 600 -450 2775 -440
rect 600 -510 605 -450
rect 660 -510 795 -450
rect 850 -510 990 -450
rect 1045 -510 1180 -450
rect 1235 -510 1375 -450
rect 1430 -510 1565 -450
rect 1620 -510 1755 -450
rect 1810 -510 1950 -450
rect 2005 -510 2140 -450
rect 2195 -510 2340 -450
rect 2765 -510 2775 -450
rect 600 -520 2775 -510
<< via2 >>
rect 130 530 460 745
rect 2340 530 2765 745
rect 130 -510 460 -450
rect 2340 -510 2765 -450
<< metal3 >>
rect -40 745 470 755
rect -40 530 130 745
rect 460 530 470 745
rect -40 -450 470 530
rect -40 -510 130 -450
rect 460 -510 470 -450
rect -40 -520 470 -510
rect 2330 745 2935 755
rect 2330 530 2340 745
rect 2765 530 2935 745
rect 2330 -450 2935 530
rect 2330 -510 2340 -450
rect 2765 -510 2935 -450
rect 2330 -520 2935 -510
use sky130_fd_pr__nfet_01v8_98DYX6  sky130_fd_pr__nfet_01v8_98DYX6_0
timestamp 1762641840
transform 1 0 1448 0 1 -410
box -1463 -310 1463 310
use sky130_fd_pr__pfet_01v8_3HM6GL  sky130_fd_pr__pfet_01v8_3HM6GL_0
timestamp 1762641840
transform 1 0 1448 0 1 469
box -1463 -519 1463 519
<< labels >>
flabel viali 1495 950 1495 950 0 FreeSans 480 0 0 0 VDD
port 3 nsew
flabel metal1 1485 -95 1485 -95 0 FreeSans 480 0 0 0 di_tg_ctrl_n
port 5 nsew
flabel viali 1495 -685 1495 -685 0 FreeSans 480 0 0 0 VSS
port 6 nsew
flabel metal1 1490 845 1490 845 0 FreeSans 480 0 0 0 di_tg_ctrl
port 8 nsew
flabel metal3 -30 -75 -30 -75 0 FreeSans 480 0 0 0 v_a
port 10 nsew
flabel metal3 2925 -75 2925 -75 0 FreeSans 480 0 0 0 v_b
port 12 nsew
<< end >>
