magic
tech sky130A
magscale 1 2
timestamp 1762641840
<< nwell >>
rect -359 -519 359 519
<< pmos >>
rect -159 -300 -129 300
rect -63 -300 -33 300
rect 33 -300 63 300
rect 129 -300 159 300
<< pdiff >>
rect -221 288 -159 300
rect -221 -288 -209 288
rect -175 -288 -159 288
rect -221 -300 -159 -288
rect -129 288 -63 300
rect -129 -288 -113 288
rect -79 -288 -63 288
rect -129 -300 -63 -288
rect -33 288 33 300
rect -33 -288 -17 288
rect 17 -288 33 288
rect -33 -300 33 -288
rect 63 288 129 300
rect 63 -288 79 288
rect 113 -288 129 288
rect 63 -300 129 -288
rect 159 288 221 300
rect 159 -288 175 288
rect 209 -288 221 288
rect 159 -300 221 -288
<< pdiffc >>
rect -209 -288 -175 288
rect -113 -288 -79 288
rect -17 -288 17 288
rect 79 -288 113 288
rect 175 -288 209 288
<< nsubdiff >>
rect -323 449 -227 483
rect 227 449 323 483
rect -323 387 -289 449
rect 289 387 323 449
rect -323 -449 -289 -387
rect 289 -449 323 -387
rect -323 -483 -227 -449
rect 227 -483 323 -449
<< nsubdiffcont >>
rect -227 449 227 483
rect -323 -387 -289 387
rect 289 -387 323 387
rect -227 -483 227 -449
<< poly >>
rect -235 395 -129 415
rect -235 360 -215 395
rect -150 360 -129 395
rect -235 340 -129 360
rect -159 300 -129 340
rect 129 395 235 415
rect 129 360 150 395
rect 215 360 235 395
rect 129 340 235 360
rect -63 300 -33 326
rect 33 300 63 326
rect 129 300 159 340
rect -159 -326 -129 -300
rect -63 -340 -33 -300
rect 33 -340 63 -300
rect 129 -326 159 -300
rect -80 -360 80 -340
rect -80 -395 -60 -360
rect 60 -395 80 -360
rect -80 -415 80 -395
<< polycont >>
rect -215 360 -150 395
rect 150 360 215 395
rect -60 -395 60 -360
<< locali >>
rect -360 505 360 520
rect -360 465 -345 505
rect 345 465 360 505
rect -360 449 -227 465
rect 227 449 360 465
rect -360 387 -289 449
rect -360 -387 -323 387
rect -235 400 -130 410
rect -235 355 -220 400
rect -175 395 -130 400
rect -150 360 -130 395
rect -175 355 -130 360
rect -235 345 -130 355
rect 130 400 235 410
rect 130 395 175 400
rect 130 360 150 395
rect 130 355 175 360
rect 220 355 235 400
rect 130 345 235 355
rect 289 387 360 449
rect -209 288 -175 304
rect -209 -304 -175 -288
rect -113 288 -79 304
rect -113 -304 -79 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 79 288 113 304
rect 79 -304 113 -288
rect 175 288 209 304
rect 175 -304 209 -288
rect -360 -449 -289 -387
rect -80 -355 80 -340
rect -80 -400 -65 -355
rect 65 -400 80 -355
rect -80 -415 80 -400
rect 323 -387 360 387
rect 289 -449 360 -387
rect -360 -483 -227 -449
rect 227 -483 360 -449
rect -360 -520 360 -483
<< viali >>
rect -345 483 345 505
rect -345 465 -227 483
rect -227 465 227 483
rect 227 465 345 483
rect -220 395 -175 400
rect -220 360 -215 395
rect -215 360 -175 395
rect -220 355 -175 360
rect 175 395 220 400
rect 175 360 215 395
rect 215 360 220 395
rect 175 355 220 360
rect -209 -288 -175 288
rect -113 -288 -79 288
rect -17 -288 17 288
rect 79 -288 113 288
rect 175 -288 209 288
rect -65 -360 65 -355
rect -65 -395 -60 -360
rect -60 -395 60 -360
rect 60 -395 65 -360
rect -65 -400 65 -395
<< metal1 >>
rect -360 505 360 520
rect -360 465 -345 505
rect 345 465 360 505
rect -360 450 360 465
rect -235 400 -160 410
rect -235 355 -220 400
rect -175 355 -160 400
rect -235 345 -160 355
rect 160 400 235 410
rect 160 355 175 400
rect 220 355 235 400
rect 160 345 235 355
rect -215 288 -169 300
rect -215 -288 -209 288
rect -175 -288 -169 288
rect -215 -300 -169 -288
rect -119 288 -73 300
rect -119 -288 -113 288
rect -79 -288 -73 288
rect -119 -300 -73 -288
rect -23 288 23 300
rect -23 -288 -17 288
rect 17 -288 23 288
rect -23 -300 23 -288
rect 73 288 119 300
rect 73 -288 79 288
rect 113 -288 119 288
rect 73 -300 119 -288
rect 169 288 215 300
rect 169 -288 175 288
rect 209 -288 215 288
rect 169 -300 215 -288
rect -80 -355 80 -340
rect -80 -400 -65 -355
rect 65 -400 80 -355
rect -80 -415 80 -400
<< labels >>
rlabel pdiffc -192 0 -192 0 0 D0
port 2 nsew
rlabel pdiffc -96 0 -96 0 0 S1
port 4 nsew
rlabel pdiffc 0 0 0 0 0 D2
port 6 nsew
rlabel pdiffc 96 0 96 0 0 S3
port 8 nsew
rlabel nsubdiffcont 0 -466 0 -466 0 B
port 1 nsew
<< properties >>
string FIXED_BBOX -306 -466 306 466
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3.0 l 0.15 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
