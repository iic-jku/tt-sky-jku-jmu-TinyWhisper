magic
tech sky130A
magscale 1 2
timestamp 1757113279
<< pwell >>
rect -11572 -782 11572 782
<< psubdiff >>
rect -11536 712 -11440 746
rect 11440 712 11536 746
rect -11536 650 -11502 712
rect 11502 650 11536 712
rect -11536 -712 -11502 -650
rect 11502 -712 11536 -650
rect -11536 -746 -11440 -712
rect 11440 -746 11536 -712
<< psubdiffcont >>
rect -11440 712 11440 746
rect -11536 -650 -11502 650
rect 11502 -650 11536 650
rect -11440 -746 11440 -712
<< xpolycontact >>
rect -11406 184 -11336 616
rect -11406 -616 -11336 -184
rect -11240 184 -11170 616
rect -11240 -616 -11170 -184
rect -11074 184 -11004 616
rect -11074 -616 -11004 -184
rect -10908 184 -10838 616
rect -10908 -616 -10838 -184
rect -10742 184 -10672 616
rect -10742 -616 -10672 -184
rect -10576 184 -10506 616
rect -10576 -616 -10506 -184
rect -10410 184 -10340 616
rect -10410 -616 -10340 -184
rect -10244 184 -10174 616
rect -10244 -616 -10174 -184
rect -10078 184 -10008 616
rect -10078 -616 -10008 -184
rect -9912 184 -9842 616
rect -9912 -616 -9842 -184
rect -9746 184 -9676 616
rect -9746 -616 -9676 -184
rect -9580 184 -9510 616
rect -9580 -616 -9510 -184
rect -9414 184 -9344 616
rect -9414 -616 -9344 -184
rect -9248 184 -9178 616
rect -9248 -616 -9178 -184
rect -9082 184 -9012 616
rect -9082 -616 -9012 -184
rect -8916 184 -8846 616
rect -8916 -616 -8846 -184
rect -8750 184 -8680 616
rect -8750 -616 -8680 -184
rect -8584 184 -8514 616
rect -8584 -616 -8514 -184
rect -8418 184 -8348 616
rect -8418 -616 -8348 -184
rect -8252 184 -8182 616
rect -8252 -616 -8182 -184
rect -8086 184 -8016 616
rect -8086 -616 -8016 -184
rect -7920 184 -7850 616
rect -7920 -616 -7850 -184
rect -7754 184 -7684 616
rect -7754 -616 -7684 -184
rect -7588 184 -7518 616
rect -7588 -616 -7518 -184
rect -7422 184 -7352 616
rect -7422 -616 -7352 -184
rect -7256 184 -7186 616
rect -7256 -616 -7186 -184
rect -7090 184 -7020 616
rect -7090 -616 -7020 -184
rect -6924 184 -6854 616
rect -6924 -616 -6854 -184
rect -6758 184 -6688 616
rect -6758 -616 -6688 -184
rect -6592 184 -6522 616
rect -6592 -616 -6522 -184
rect -6426 184 -6356 616
rect -6426 -616 -6356 -184
rect -6260 184 -6190 616
rect -6260 -616 -6190 -184
rect -6094 184 -6024 616
rect -6094 -616 -6024 -184
rect -5928 184 -5858 616
rect -5928 -616 -5858 -184
rect -5762 184 -5692 616
rect -5762 -616 -5692 -184
rect -5596 184 -5526 616
rect -5596 -616 -5526 -184
rect -5430 184 -5360 616
rect -5430 -616 -5360 -184
rect -5264 184 -5194 616
rect -5264 -616 -5194 -184
rect -5098 184 -5028 616
rect -5098 -616 -5028 -184
rect -4932 184 -4862 616
rect -4932 -616 -4862 -184
rect -4766 184 -4696 616
rect -4766 -616 -4696 -184
rect -4600 184 -4530 616
rect -4600 -616 -4530 -184
rect -4434 184 -4364 616
rect -4434 -616 -4364 -184
rect -4268 184 -4198 616
rect -4268 -616 -4198 -184
rect -4102 184 -4032 616
rect -4102 -616 -4032 -184
rect -3936 184 -3866 616
rect -3936 -616 -3866 -184
rect -3770 184 -3700 616
rect -3770 -616 -3700 -184
rect -3604 184 -3534 616
rect -3604 -616 -3534 -184
rect -3438 184 -3368 616
rect -3438 -616 -3368 -184
rect -3272 184 -3202 616
rect -3272 -616 -3202 -184
rect -3106 184 -3036 616
rect -3106 -616 -3036 -184
rect -2940 184 -2870 616
rect -2940 -616 -2870 -184
rect -2774 184 -2704 616
rect -2774 -616 -2704 -184
rect -2608 184 -2538 616
rect -2608 -616 -2538 -184
rect -2442 184 -2372 616
rect -2442 -616 -2372 -184
rect -2276 184 -2206 616
rect -2276 -616 -2206 -184
rect -2110 184 -2040 616
rect -2110 -616 -2040 -184
rect -1944 184 -1874 616
rect -1944 -616 -1874 -184
rect -1778 184 -1708 616
rect -1778 -616 -1708 -184
rect -1612 184 -1542 616
rect -1612 -616 -1542 -184
rect -1446 184 -1376 616
rect -1446 -616 -1376 -184
rect -1280 184 -1210 616
rect -1280 -616 -1210 -184
rect -1114 184 -1044 616
rect -1114 -616 -1044 -184
rect -948 184 -878 616
rect -948 -616 -878 -184
rect -782 184 -712 616
rect -782 -616 -712 -184
rect -616 184 -546 616
rect -616 -616 -546 -184
rect -450 184 -380 616
rect -450 -616 -380 -184
rect -284 184 -214 616
rect -284 -616 -214 -184
rect -118 184 -48 616
rect -118 -616 -48 -184
rect 48 184 118 616
rect 48 -616 118 -184
rect 214 184 284 616
rect 214 -616 284 -184
rect 380 184 450 616
rect 380 -616 450 -184
rect 546 184 616 616
rect 546 -616 616 -184
rect 712 184 782 616
rect 712 -616 782 -184
rect 878 184 948 616
rect 878 -616 948 -184
rect 1044 184 1114 616
rect 1044 -616 1114 -184
rect 1210 184 1280 616
rect 1210 -616 1280 -184
rect 1376 184 1446 616
rect 1376 -616 1446 -184
rect 1542 184 1612 616
rect 1542 -616 1612 -184
rect 1708 184 1778 616
rect 1708 -616 1778 -184
rect 1874 184 1944 616
rect 1874 -616 1944 -184
rect 2040 184 2110 616
rect 2040 -616 2110 -184
rect 2206 184 2276 616
rect 2206 -616 2276 -184
rect 2372 184 2442 616
rect 2372 -616 2442 -184
rect 2538 184 2608 616
rect 2538 -616 2608 -184
rect 2704 184 2774 616
rect 2704 -616 2774 -184
rect 2870 184 2940 616
rect 2870 -616 2940 -184
rect 3036 184 3106 616
rect 3036 -616 3106 -184
rect 3202 184 3272 616
rect 3202 -616 3272 -184
rect 3368 184 3438 616
rect 3368 -616 3438 -184
rect 3534 184 3604 616
rect 3534 -616 3604 -184
rect 3700 184 3770 616
rect 3700 -616 3770 -184
rect 3866 184 3936 616
rect 3866 -616 3936 -184
rect 4032 184 4102 616
rect 4032 -616 4102 -184
rect 4198 184 4268 616
rect 4198 -616 4268 -184
rect 4364 184 4434 616
rect 4364 -616 4434 -184
rect 4530 184 4600 616
rect 4530 -616 4600 -184
rect 4696 184 4766 616
rect 4696 -616 4766 -184
rect 4862 184 4932 616
rect 4862 -616 4932 -184
rect 5028 184 5098 616
rect 5028 -616 5098 -184
rect 5194 184 5264 616
rect 5194 -616 5264 -184
rect 5360 184 5430 616
rect 5360 -616 5430 -184
rect 5526 184 5596 616
rect 5526 -616 5596 -184
rect 5692 184 5762 616
rect 5692 -616 5762 -184
rect 5858 184 5928 616
rect 5858 -616 5928 -184
rect 6024 184 6094 616
rect 6024 -616 6094 -184
rect 6190 184 6260 616
rect 6190 -616 6260 -184
rect 6356 184 6426 616
rect 6356 -616 6426 -184
rect 6522 184 6592 616
rect 6522 -616 6592 -184
rect 6688 184 6758 616
rect 6688 -616 6758 -184
rect 6854 184 6924 616
rect 6854 -616 6924 -184
rect 7020 184 7090 616
rect 7020 -616 7090 -184
rect 7186 184 7256 616
rect 7186 -616 7256 -184
rect 7352 184 7422 616
rect 7352 -616 7422 -184
rect 7518 184 7588 616
rect 7518 -616 7588 -184
rect 7684 184 7754 616
rect 7684 -616 7754 -184
rect 7850 184 7920 616
rect 7850 -616 7920 -184
rect 8016 184 8086 616
rect 8016 -616 8086 -184
rect 8182 184 8252 616
rect 8182 -616 8252 -184
rect 8348 184 8418 616
rect 8348 -616 8418 -184
rect 8514 184 8584 616
rect 8514 -616 8584 -184
rect 8680 184 8750 616
rect 8680 -616 8750 -184
rect 8846 184 8916 616
rect 8846 -616 8916 -184
rect 9012 184 9082 616
rect 9012 -616 9082 -184
rect 9178 184 9248 616
rect 9178 -616 9248 -184
rect 9344 184 9414 616
rect 9344 -616 9414 -184
rect 9510 184 9580 616
rect 9510 -616 9580 -184
rect 9676 184 9746 616
rect 9676 -616 9746 -184
rect 9842 184 9912 616
rect 9842 -616 9912 -184
rect 10008 184 10078 616
rect 10008 -616 10078 -184
rect 10174 184 10244 616
rect 10174 -616 10244 -184
rect 10340 184 10410 616
rect 10340 -616 10410 -184
rect 10506 184 10576 616
rect 10506 -616 10576 -184
rect 10672 184 10742 616
rect 10672 -616 10742 -184
rect 10838 184 10908 616
rect 10838 -616 10908 -184
rect 11004 184 11074 616
rect 11004 -616 11074 -184
rect 11170 184 11240 616
rect 11170 -616 11240 -184
rect 11336 184 11406 616
rect 11336 -616 11406 -184
<< xpolyres >>
rect -11406 -184 -11336 184
rect -11240 -184 -11170 184
rect -11074 -184 -11004 184
rect -10908 -184 -10838 184
rect -10742 -184 -10672 184
rect -10576 -184 -10506 184
rect -10410 -184 -10340 184
rect -10244 -184 -10174 184
rect -10078 -184 -10008 184
rect -9912 -184 -9842 184
rect -9746 -184 -9676 184
rect -9580 -184 -9510 184
rect -9414 -184 -9344 184
rect -9248 -184 -9178 184
rect -9082 -184 -9012 184
rect -8916 -184 -8846 184
rect -8750 -184 -8680 184
rect -8584 -184 -8514 184
rect -8418 -184 -8348 184
rect -8252 -184 -8182 184
rect -8086 -184 -8016 184
rect -7920 -184 -7850 184
rect -7754 -184 -7684 184
rect -7588 -184 -7518 184
rect -7422 -184 -7352 184
rect -7256 -184 -7186 184
rect -7090 -184 -7020 184
rect -6924 -184 -6854 184
rect -6758 -184 -6688 184
rect -6592 -184 -6522 184
rect -6426 -184 -6356 184
rect -6260 -184 -6190 184
rect -6094 -184 -6024 184
rect -5928 -184 -5858 184
rect -5762 -184 -5692 184
rect -5596 -184 -5526 184
rect -5430 -184 -5360 184
rect -5264 -184 -5194 184
rect -5098 -184 -5028 184
rect -4932 -184 -4862 184
rect -4766 -184 -4696 184
rect -4600 -184 -4530 184
rect -4434 -184 -4364 184
rect -4268 -184 -4198 184
rect -4102 -184 -4032 184
rect -3936 -184 -3866 184
rect -3770 -184 -3700 184
rect -3604 -184 -3534 184
rect -3438 -184 -3368 184
rect -3272 -184 -3202 184
rect -3106 -184 -3036 184
rect -2940 -184 -2870 184
rect -2774 -184 -2704 184
rect -2608 -184 -2538 184
rect -2442 -184 -2372 184
rect -2276 -184 -2206 184
rect -2110 -184 -2040 184
rect -1944 -184 -1874 184
rect -1778 -184 -1708 184
rect -1612 -184 -1542 184
rect -1446 -184 -1376 184
rect -1280 -184 -1210 184
rect -1114 -184 -1044 184
rect -948 -184 -878 184
rect -782 -184 -712 184
rect -616 -184 -546 184
rect -450 -184 -380 184
rect -284 -184 -214 184
rect -118 -184 -48 184
rect 48 -184 118 184
rect 214 -184 284 184
rect 380 -184 450 184
rect 546 -184 616 184
rect 712 -184 782 184
rect 878 -184 948 184
rect 1044 -184 1114 184
rect 1210 -184 1280 184
rect 1376 -184 1446 184
rect 1542 -184 1612 184
rect 1708 -184 1778 184
rect 1874 -184 1944 184
rect 2040 -184 2110 184
rect 2206 -184 2276 184
rect 2372 -184 2442 184
rect 2538 -184 2608 184
rect 2704 -184 2774 184
rect 2870 -184 2940 184
rect 3036 -184 3106 184
rect 3202 -184 3272 184
rect 3368 -184 3438 184
rect 3534 -184 3604 184
rect 3700 -184 3770 184
rect 3866 -184 3936 184
rect 4032 -184 4102 184
rect 4198 -184 4268 184
rect 4364 -184 4434 184
rect 4530 -184 4600 184
rect 4696 -184 4766 184
rect 4862 -184 4932 184
rect 5028 -184 5098 184
rect 5194 -184 5264 184
rect 5360 -184 5430 184
rect 5526 -184 5596 184
rect 5692 -184 5762 184
rect 5858 -184 5928 184
rect 6024 -184 6094 184
rect 6190 -184 6260 184
rect 6356 -184 6426 184
rect 6522 -184 6592 184
rect 6688 -184 6758 184
rect 6854 -184 6924 184
rect 7020 -184 7090 184
rect 7186 -184 7256 184
rect 7352 -184 7422 184
rect 7518 -184 7588 184
rect 7684 -184 7754 184
rect 7850 -184 7920 184
rect 8016 -184 8086 184
rect 8182 -184 8252 184
rect 8348 -184 8418 184
rect 8514 -184 8584 184
rect 8680 -184 8750 184
rect 8846 -184 8916 184
rect 9012 -184 9082 184
rect 9178 -184 9248 184
rect 9344 -184 9414 184
rect 9510 -184 9580 184
rect 9676 -184 9746 184
rect 9842 -184 9912 184
rect 10008 -184 10078 184
rect 10174 -184 10244 184
rect 10340 -184 10410 184
rect 10506 -184 10576 184
rect 10672 -184 10742 184
rect 10838 -184 10908 184
rect 11004 -184 11074 184
rect 11170 -184 11240 184
rect 11336 -184 11406 184
<< locali >>
rect -11536 712 -11440 746
rect 11440 712 11536 746
rect -11536 650 -11502 712
rect 11502 650 11536 712
rect -11536 -712 -11502 -650
rect 11502 -712 11536 -650
rect -11536 -746 -11440 -712
rect 11440 -746 11536 -712
<< viali >>
rect -11390 201 -11352 598
rect -11224 201 -11186 598
rect -11058 201 -11020 598
rect -10892 201 -10854 598
rect -10726 201 -10688 598
rect -10560 201 -10522 598
rect -10394 201 -10356 598
rect -10228 201 -10190 598
rect -10062 201 -10024 598
rect -9896 201 -9858 598
rect -9730 201 -9692 598
rect -9564 201 -9526 598
rect -9398 201 -9360 598
rect -9232 201 -9194 598
rect -9066 201 -9028 598
rect -8900 201 -8862 598
rect -8734 201 -8696 598
rect -8568 201 -8530 598
rect -8402 201 -8364 598
rect -8236 201 -8198 598
rect -8070 201 -8032 598
rect -7904 201 -7866 598
rect -7738 201 -7700 598
rect -7572 201 -7534 598
rect -7406 201 -7368 598
rect -7240 201 -7202 598
rect -7074 201 -7036 598
rect -6908 201 -6870 598
rect -6742 201 -6704 598
rect -6576 201 -6538 598
rect -6410 201 -6372 598
rect -6244 201 -6206 598
rect -6078 201 -6040 598
rect -5912 201 -5874 598
rect -5746 201 -5708 598
rect -5580 201 -5542 598
rect -5414 201 -5376 598
rect -5248 201 -5210 598
rect -5082 201 -5044 598
rect -4916 201 -4878 598
rect -4750 201 -4712 598
rect -4584 201 -4546 598
rect -4418 201 -4380 598
rect -4252 201 -4214 598
rect -4086 201 -4048 598
rect -3920 201 -3882 598
rect -3754 201 -3716 598
rect -3588 201 -3550 598
rect -3422 201 -3384 598
rect -3256 201 -3218 598
rect -3090 201 -3052 598
rect -2924 201 -2886 598
rect -2758 201 -2720 598
rect -2592 201 -2554 598
rect -2426 201 -2388 598
rect -2260 201 -2222 598
rect -2094 201 -2056 598
rect -1928 201 -1890 598
rect -1762 201 -1724 598
rect -1596 201 -1558 598
rect -1430 201 -1392 598
rect -1264 201 -1226 598
rect -1098 201 -1060 598
rect -932 201 -894 598
rect -766 201 -728 598
rect -600 201 -562 598
rect -434 201 -396 598
rect -268 201 -230 598
rect -102 201 -64 598
rect 64 201 102 598
rect 230 201 268 598
rect 396 201 434 598
rect 562 201 600 598
rect 728 201 766 598
rect 894 201 932 598
rect 1060 201 1098 598
rect 1226 201 1264 598
rect 1392 201 1430 598
rect 1558 201 1596 598
rect 1724 201 1762 598
rect 1890 201 1928 598
rect 2056 201 2094 598
rect 2222 201 2260 598
rect 2388 201 2426 598
rect 2554 201 2592 598
rect 2720 201 2758 598
rect 2886 201 2924 598
rect 3052 201 3090 598
rect 3218 201 3256 598
rect 3384 201 3422 598
rect 3550 201 3588 598
rect 3716 201 3754 598
rect 3882 201 3920 598
rect 4048 201 4086 598
rect 4214 201 4252 598
rect 4380 201 4418 598
rect 4546 201 4584 598
rect 4712 201 4750 598
rect 4878 201 4916 598
rect 5044 201 5082 598
rect 5210 201 5248 598
rect 5376 201 5414 598
rect 5542 201 5580 598
rect 5708 201 5746 598
rect 5874 201 5912 598
rect 6040 201 6078 598
rect 6206 201 6244 598
rect 6372 201 6410 598
rect 6538 201 6576 598
rect 6704 201 6742 598
rect 6870 201 6908 598
rect 7036 201 7074 598
rect 7202 201 7240 598
rect 7368 201 7406 598
rect 7534 201 7572 598
rect 7700 201 7738 598
rect 7866 201 7904 598
rect 8032 201 8070 598
rect 8198 201 8236 598
rect 8364 201 8402 598
rect 8530 201 8568 598
rect 8696 201 8734 598
rect 8862 201 8900 598
rect 9028 201 9066 598
rect 9194 201 9232 598
rect 9360 201 9398 598
rect 9526 201 9564 598
rect 9692 201 9730 598
rect 9858 201 9896 598
rect 10024 201 10062 598
rect 10190 201 10228 598
rect 10356 201 10394 598
rect 10522 201 10560 598
rect 10688 201 10726 598
rect 10854 201 10892 598
rect 11020 201 11058 598
rect 11186 201 11224 598
rect 11352 201 11390 598
rect -11390 -598 -11352 -201
rect -11224 -598 -11186 -201
rect -11058 -598 -11020 -201
rect -10892 -598 -10854 -201
rect -10726 -598 -10688 -201
rect -10560 -598 -10522 -201
rect -10394 -598 -10356 -201
rect -10228 -598 -10190 -201
rect -10062 -598 -10024 -201
rect -9896 -598 -9858 -201
rect -9730 -598 -9692 -201
rect -9564 -598 -9526 -201
rect -9398 -598 -9360 -201
rect -9232 -598 -9194 -201
rect -9066 -598 -9028 -201
rect -8900 -598 -8862 -201
rect -8734 -598 -8696 -201
rect -8568 -598 -8530 -201
rect -8402 -598 -8364 -201
rect -8236 -598 -8198 -201
rect -8070 -598 -8032 -201
rect -7904 -598 -7866 -201
rect -7738 -598 -7700 -201
rect -7572 -598 -7534 -201
rect -7406 -598 -7368 -201
rect -7240 -598 -7202 -201
rect -7074 -598 -7036 -201
rect -6908 -598 -6870 -201
rect -6742 -598 -6704 -201
rect -6576 -598 -6538 -201
rect -6410 -598 -6372 -201
rect -6244 -598 -6206 -201
rect -6078 -598 -6040 -201
rect -5912 -598 -5874 -201
rect -5746 -598 -5708 -201
rect -5580 -598 -5542 -201
rect -5414 -598 -5376 -201
rect -5248 -598 -5210 -201
rect -5082 -598 -5044 -201
rect -4916 -598 -4878 -201
rect -4750 -598 -4712 -201
rect -4584 -598 -4546 -201
rect -4418 -598 -4380 -201
rect -4252 -598 -4214 -201
rect -4086 -598 -4048 -201
rect -3920 -598 -3882 -201
rect -3754 -598 -3716 -201
rect -3588 -598 -3550 -201
rect -3422 -598 -3384 -201
rect -3256 -598 -3218 -201
rect -3090 -598 -3052 -201
rect -2924 -598 -2886 -201
rect -2758 -598 -2720 -201
rect -2592 -598 -2554 -201
rect -2426 -598 -2388 -201
rect -2260 -598 -2222 -201
rect -2094 -598 -2056 -201
rect -1928 -598 -1890 -201
rect -1762 -598 -1724 -201
rect -1596 -598 -1558 -201
rect -1430 -598 -1392 -201
rect -1264 -598 -1226 -201
rect -1098 -598 -1060 -201
rect -932 -598 -894 -201
rect -766 -598 -728 -201
rect -600 -598 -562 -201
rect -434 -598 -396 -201
rect -268 -598 -230 -201
rect -102 -598 -64 -201
rect 64 -598 102 -201
rect 230 -598 268 -201
rect 396 -598 434 -201
rect 562 -598 600 -201
rect 728 -598 766 -201
rect 894 -598 932 -201
rect 1060 -598 1098 -201
rect 1226 -598 1264 -201
rect 1392 -598 1430 -201
rect 1558 -598 1596 -201
rect 1724 -598 1762 -201
rect 1890 -598 1928 -201
rect 2056 -598 2094 -201
rect 2222 -598 2260 -201
rect 2388 -598 2426 -201
rect 2554 -598 2592 -201
rect 2720 -598 2758 -201
rect 2886 -598 2924 -201
rect 3052 -598 3090 -201
rect 3218 -598 3256 -201
rect 3384 -598 3422 -201
rect 3550 -598 3588 -201
rect 3716 -598 3754 -201
rect 3882 -598 3920 -201
rect 4048 -598 4086 -201
rect 4214 -598 4252 -201
rect 4380 -598 4418 -201
rect 4546 -598 4584 -201
rect 4712 -598 4750 -201
rect 4878 -598 4916 -201
rect 5044 -598 5082 -201
rect 5210 -598 5248 -201
rect 5376 -598 5414 -201
rect 5542 -598 5580 -201
rect 5708 -598 5746 -201
rect 5874 -598 5912 -201
rect 6040 -598 6078 -201
rect 6206 -598 6244 -201
rect 6372 -598 6410 -201
rect 6538 -598 6576 -201
rect 6704 -598 6742 -201
rect 6870 -598 6908 -201
rect 7036 -598 7074 -201
rect 7202 -598 7240 -201
rect 7368 -598 7406 -201
rect 7534 -598 7572 -201
rect 7700 -598 7738 -201
rect 7866 -598 7904 -201
rect 8032 -598 8070 -201
rect 8198 -598 8236 -201
rect 8364 -598 8402 -201
rect 8530 -598 8568 -201
rect 8696 -598 8734 -201
rect 8862 -598 8900 -201
rect 9028 -598 9066 -201
rect 9194 -598 9232 -201
rect 9360 -598 9398 -201
rect 9526 -598 9564 -201
rect 9692 -598 9730 -201
rect 9858 -598 9896 -201
rect 10024 -598 10062 -201
rect 10190 -598 10228 -201
rect 10356 -598 10394 -201
rect 10522 -598 10560 -201
rect 10688 -598 10726 -201
rect 10854 -598 10892 -201
rect 11020 -598 11058 -201
rect 11186 -598 11224 -201
rect 11352 -598 11390 -201
<< metal1 >>
rect -11396 598 -11346 610
rect -11396 201 -11390 598
rect -11352 201 -11346 598
rect -11396 189 -11346 201
rect -11230 598 -11180 610
rect -11230 201 -11224 598
rect -11186 201 -11180 598
rect -11230 189 -11180 201
rect -11064 598 -11014 610
rect -11064 201 -11058 598
rect -11020 201 -11014 598
rect -11064 189 -11014 201
rect -10898 598 -10848 610
rect -10898 201 -10892 598
rect -10854 201 -10848 598
rect -10898 189 -10848 201
rect -10732 598 -10682 610
rect -10732 201 -10726 598
rect -10688 201 -10682 598
rect -10732 189 -10682 201
rect -10566 598 -10516 610
rect -10566 201 -10560 598
rect -10522 201 -10516 598
rect -10566 189 -10516 201
rect -10400 598 -10350 610
rect -10400 201 -10394 598
rect -10356 201 -10350 598
rect -10400 189 -10350 201
rect -10234 598 -10184 610
rect -10234 201 -10228 598
rect -10190 201 -10184 598
rect -10234 189 -10184 201
rect -10068 598 -10018 610
rect -10068 201 -10062 598
rect -10024 201 -10018 598
rect -10068 189 -10018 201
rect -9902 598 -9852 610
rect -9902 201 -9896 598
rect -9858 201 -9852 598
rect -9902 189 -9852 201
rect -9736 598 -9686 610
rect -9736 201 -9730 598
rect -9692 201 -9686 598
rect -9736 189 -9686 201
rect -9570 598 -9520 610
rect -9570 201 -9564 598
rect -9526 201 -9520 598
rect -9570 189 -9520 201
rect -9404 598 -9354 610
rect -9404 201 -9398 598
rect -9360 201 -9354 598
rect -9404 189 -9354 201
rect -9238 598 -9188 610
rect -9238 201 -9232 598
rect -9194 201 -9188 598
rect -9238 189 -9188 201
rect -9072 598 -9022 610
rect -9072 201 -9066 598
rect -9028 201 -9022 598
rect -9072 189 -9022 201
rect -8906 598 -8856 610
rect -8906 201 -8900 598
rect -8862 201 -8856 598
rect -8906 189 -8856 201
rect -8740 598 -8690 610
rect -8740 201 -8734 598
rect -8696 201 -8690 598
rect -8740 189 -8690 201
rect -8574 598 -8524 610
rect -8574 201 -8568 598
rect -8530 201 -8524 598
rect -8574 189 -8524 201
rect -8408 598 -8358 610
rect -8408 201 -8402 598
rect -8364 201 -8358 598
rect -8408 189 -8358 201
rect -8242 598 -8192 610
rect -8242 201 -8236 598
rect -8198 201 -8192 598
rect -8242 189 -8192 201
rect -8076 598 -8026 610
rect -8076 201 -8070 598
rect -8032 201 -8026 598
rect -8076 189 -8026 201
rect -7910 598 -7860 610
rect -7910 201 -7904 598
rect -7866 201 -7860 598
rect -7910 189 -7860 201
rect -7744 598 -7694 610
rect -7744 201 -7738 598
rect -7700 201 -7694 598
rect -7744 189 -7694 201
rect -7578 598 -7528 610
rect -7578 201 -7572 598
rect -7534 201 -7528 598
rect -7578 189 -7528 201
rect -7412 598 -7362 610
rect -7412 201 -7406 598
rect -7368 201 -7362 598
rect -7412 189 -7362 201
rect -7246 598 -7196 610
rect -7246 201 -7240 598
rect -7202 201 -7196 598
rect -7246 189 -7196 201
rect -7080 598 -7030 610
rect -7080 201 -7074 598
rect -7036 201 -7030 598
rect -7080 189 -7030 201
rect -6914 598 -6864 610
rect -6914 201 -6908 598
rect -6870 201 -6864 598
rect -6914 189 -6864 201
rect -6748 598 -6698 610
rect -6748 201 -6742 598
rect -6704 201 -6698 598
rect -6748 189 -6698 201
rect -6582 598 -6532 610
rect -6582 201 -6576 598
rect -6538 201 -6532 598
rect -6582 189 -6532 201
rect -6416 598 -6366 610
rect -6416 201 -6410 598
rect -6372 201 -6366 598
rect -6416 189 -6366 201
rect -6250 598 -6200 610
rect -6250 201 -6244 598
rect -6206 201 -6200 598
rect -6250 189 -6200 201
rect -6084 598 -6034 610
rect -6084 201 -6078 598
rect -6040 201 -6034 598
rect -6084 189 -6034 201
rect -5918 598 -5868 610
rect -5918 201 -5912 598
rect -5874 201 -5868 598
rect -5918 189 -5868 201
rect -5752 598 -5702 610
rect -5752 201 -5746 598
rect -5708 201 -5702 598
rect -5752 189 -5702 201
rect -5586 598 -5536 610
rect -5586 201 -5580 598
rect -5542 201 -5536 598
rect -5586 189 -5536 201
rect -5420 598 -5370 610
rect -5420 201 -5414 598
rect -5376 201 -5370 598
rect -5420 189 -5370 201
rect -5254 598 -5204 610
rect -5254 201 -5248 598
rect -5210 201 -5204 598
rect -5254 189 -5204 201
rect -5088 598 -5038 610
rect -5088 201 -5082 598
rect -5044 201 -5038 598
rect -5088 189 -5038 201
rect -4922 598 -4872 610
rect -4922 201 -4916 598
rect -4878 201 -4872 598
rect -4922 189 -4872 201
rect -4756 598 -4706 610
rect -4756 201 -4750 598
rect -4712 201 -4706 598
rect -4756 189 -4706 201
rect -4590 598 -4540 610
rect -4590 201 -4584 598
rect -4546 201 -4540 598
rect -4590 189 -4540 201
rect -4424 598 -4374 610
rect -4424 201 -4418 598
rect -4380 201 -4374 598
rect -4424 189 -4374 201
rect -4258 598 -4208 610
rect -4258 201 -4252 598
rect -4214 201 -4208 598
rect -4258 189 -4208 201
rect -4092 598 -4042 610
rect -4092 201 -4086 598
rect -4048 201 -4042 598
rect -4092 189 -4042 201
rect -3926 598 -3876 610
rect -3926 201 -3920 598
rect -3882 201 -3876 598
rect -3926 189 -3876 201
rect -3760 598 -3710 610
rect -3760 201 -3754 598
rect -3716 201 -3710 598
rect -3760 189 -3710 201
rect -3594 598 -3544 610
rect -3594 201 -3588 598
rect -3550 201 -3544 598
rect -3594 189 -3544 201
rect -3428 598 -3378 610
rect -3428 201 -3422 598
rect -3384 201 -3378 598
rect -3428 189 -3378 201
rect -3262 598 -3212 610
rect -3262 201 -3256 598
rect -3218 201 -3212 598
rect -3262 189 -3212 201
rect -3096 598 -3046 610
rect -3096 201 -3090 598
rect -3052 201 -3046 598
rect -3096 189 -3046 201
rect -2930 598 -2880 610
rect -2930 201 -2924 598
rect -2886 201 -2880 598
rect -2930 189 -2880 201
rect -2764 598 -2714 610
rect -2764 201 -2758 598
rect -2720 201 -2714 598
rect -2764 189 -2714 201
rect -2598 598 -2548 610
rect -2598 201 -2592 598
rect -2554 201 -2548 598
rect -2598 189 -2548 201
rect -2432 598 -2382 610
rect -2432 201 -2426 598
rect -2388 201 -2382 598
rect -2432 189 -2382 201
rect -2266 598 -2216 610
rect -2266 201 -2260 598
rect -2222 201 -2216 598
rect -2266 189 -2216 201
rect -2100 598 -2050 610
rect -2100 201 -2094 598
rect -2056 201 -2050 598
rect -2100 189 -2050 201
rect -1934 598 -1884 610
rect -1934 201 -1928 598
rect -1890 201 -1884 598
rect -1934 189 -1884 201
rect -1768 598 -1718 610
rect -1768 201 -1762 598
rect -1724 201 -1718 598
rect -1768 189 -1718 201
rect -1602 598 -1552 610
rect -1602 201 -1596 598
rect -1558 201 -1552 598
rect -1602 189 -1552 201
rect -1436 598 -1386 610
rect -1436 201 -1430 598
rect -1392 201 -1386 598
rect -1436 189 -1386 201
rect -1270 598 -1220 610
rect -1270 201 -1264 598
rect -1226 201 -1220 598
rect -1270 189 -1220 201
rect -1104 598 -1054 610
rect -1104 201 -1098 598
rect -1060 201 -1054 598
rect -1104 189 -1054 201
rect -938 598 -888 610
rect -938 201 -932 598
rect -894 201 -888 598
rect -938 189 -888 201
rect -772 598 -722 610
rect -772 201 -766 598
rect -728 201 -722 598
rect -772 189 -722 201
rect -606 598 -556 610
rect -606 201 -600 598
rect -562 201 -556 598
rect -606 189 -556 201
rect -440 598 -390 610
rect -440 201 -434 598
rect -396 201 -390 598
rect -440 189 -390 201
rect -274 598 -224 610
rect -274 201 -268 598
rect -230 201 -224 598
rect -274 189 -224 201
rect -108 598 -58 610
rect -108 201 -102 598
rect -64 201 -58 598
rect -108 189 -58 201
rect 58 598 108 610
rect 58 201 64 598
rect 102 201 108 598
rect 58 189 108 201
rect 224 598 274 610
rect 224 201 230 598
rect 268 201 274 598
rect 224 189 274 201
rect 390 598 440 610
rect 390 201 396 598
rect 434 201 440 598
rect 390 189 440 201
rect 556 598 606 610
rect 556 201 562 598
rect 600 201 606 598
rect 556 189 606 201
rect 722 598 772 610
rect 722 201 728 598
rect 766 201 772 598
rect 722 189 772 201
rect 888 598 938 610
rect 888 201 894 598
rect 932 201 938 598
rect 888 189 938 201
rect 1054 598 1104 610
rect 1054 201 1060 598
rect 1098 201 1104 598
rect 1054 189 1104 201
rect 1220 598 1270 610
rect 1220 201 1226 598
rect 1264 201 1270 598
rect 1220 189 1270 201
rect 1386 598 1436 610
rect 1386 201 1392 598
rect 1430 201 1436 598
rect 1386 189 1436 201
rect 1552 598 1602 610
rect 1552 201 1558 598
rect 1596 201 1602 598
rect 1552 189 1602 201
rect 1718 598 1768 610
rect 1718 201 1724 598
rect 1762 201 1768 598
rect 1718 189 1768 201
rect 1884 598 1934 610
rect 1884 201 1890 598
rect 1928 201 1934 598
rect 1884 189 1934 201
rect 2050 598 2100 610
rect 2050 201 2056 598
rect 2094 201 2100 598
rect 2050 189 2100 201
rect 2216 598 2266 610
rect 2216 201 2222 598
rect 2260 201 2266 598
rect 2216 189 2266 201
rect 2382 598 2432 610
rect 2382 201 2388 598
rect 2426 201 2432 598
rect 2382 189 2432 201
rect 2548 598 2598 610
rect 2548 201 2554 598
rect 2592 201 2598 598
rect 2548 189 2598 201
rect 2714 598 2764 610
rect 2714 201 2720 598
rect 2758 201 2764 598
rect 2714 189 2764 201
rect 2880 598 2930 610
rect 2880 201 2886 598
rect 2924 201 2930 598
rect 2880 189 2930 201
rect 3046 598 3096 610
rect 3046 201 3052 598
rect 3090 201 3096 598
rect 3046 189 3096 201
rect 3212 598 3262 610
rect 3212 201 3218 598
rect 3256 201 3262 598
rect 3212 189 3262 201
rect 3378 598 3428 610
rect 3378 201 3384 598
rect 3422 201 3428 598
rect 3378 189 3428 201
rect 3544 598 3594 610
rect 3544 201 3550 598
rect 3588 201 3594 598
rect 3544 189 3594 201
rect 3710 598 3760 610
rect 3710 201 3716 598
rect 3754 201 3760 598
rect 3710 189 3760 201
rect 3876 598 3926 610
rect 3876 201 3882 598
rect 3920 201 3926 598
rect 3876 189 3926 201
rect 4042 598 4092 610
rect 4042 201 4048 598
rect 4086 201 4092 598
rect 4042 189 4092 201
rect 4208 598 4258 610
rect 4208 201 4214 598
rect 4252 201 4258 598
rect 4208 189 4258 201
rect 4374 598 4424 610
rect 4374 201 4380 598
rect 4418 201 4424 598
rect 4374 189 4424 201
rect 4540 598 4590 610
rect 4540 201 4546 598
rect 4584 201 4590 598
rect 4540 189 4590 201
rect 4706 598 4756 610
rect 4706 201 4712 598
rect 4750 201 4756 598
rect 4706 189 4756 201
rect 4872 598 4922 610
rect 4872 201 4878 598
rect 4916 201 4922 598
rect 4872 189 4922 201
rect 5038 598 5088 610
rect 5038 201 5044 598
rect 5082 201 5088 598
rect 5038 189 5088 201
rect 5204 598 5254 610
rect 5204 201 5210 598
rect 5248 201 5254 598
rect 5204 189 5254 201
rect 5370 598 5420 610
rect 5370 201 5376 598
rect 5414 201 5420 598
rect 5370 189 5420 201
rect 5536 598 5586 610
rect 5536 201 5542 598
rect 5580 201 5586 598
rect 5536 189 5586 201
rect 5702 598 5752 610
rect 5702 201 5708 598
rect 5746 201 5752 598
rect 5702 189 5752 201
rect 5868 598 5918 610
rect 5868 201 5874 598
rect 5912 201 5918 598
rect 5868 189 5918 201
rect 6034 598 6084 610
rect 6034 201 6040 598
rect 6078 201 6084 598
rect 6034 189 6084 201
rect 6200 598 6250 610
rect 6200 201 6206 598
rect 6244 201 6250 598
rect 6200 189 6250 201
rect 6366 598 6416 610
rect 6366 201 6372 598
rect 6410 201 6416 598
rect 6366 189 6416 201
rect 6532 598 6582 610
rect 6532 201 6538 598
rect 6576 201 6582 598
rect 6532 189 6582 201
rect 6698 598 6748 610
rect 6698 201 6704 598
rect 6742 201 6748 598
rect 6698 189 6748 201
rect 6864 598 6914 610
rect 6864 201 6870 598
rect 6908 201 6914 598
rect 6864 189 6914 201
rect 7030 598 7080 610
rect 7030 201 7036 598
rect 7074 201 7080 598
rect 7030 189 7080 201
rect 7196 598 7246 610
rect 7196 201 7202 598
rect 7240 201 7246 598
rect 7196 189 7246 201
rect 7362 598 7412 610
rect 7362 201 7368 598
rect 7406 201 7412 598
rect 7362 189 7412 201
rect 7528 598 7578 610
rect 7528 201 7534 598
rect 7572 201 7578 598
rect 7528 189 7578 201
rect 7694 598 7744 610
rect 7694 201 7700 598
rect 7738 201 7744 598
rect 7694 189 7744 201
rect 7860 598 7910 610
rect 7860 201 7866 598
rect 7904 201 7910 598
rect 7860 189 7910 201
rect 8026 598 8076 610
rect 8026 201 8032 598
rect 8070 201 8076 598
rect 8026 189 8076 201
rect 8192 598 8242 610
rect 8192 201 8198 598
rect 8236 201 8242 598
rect 8192 189 8242 201
rect 8358 598 8408 610
rect 8358 201 8364 598
rect 8402 201 8408 598
rect 8358 189 8408 201
rect 8524 598 8574 610
rect 8524 201 8530 598
rect 8568 201 8574 598
rect 8524 189 8574 201
rect 8690 598 8740 610
rect 8690 201 8696 598
rect 8734 201 8740 598
rect 8690 189 8740 201
rect 8856 598 8906 610
rect 8856 201 8862 598
rect 8900 201 8906 598
rect 8856 189 8906 201
rect 9022 598 9072 610
rect 9022 201 9028 598
rect 9066 201 9072 598
rect 9022 189 9072 201
rect 9188 598 9238 610
rect 9188 201 9194 598
rect 9232 201 9238 598
rect 9188 189 9238 201
rect 9354 598 9404 610
rect 9354 201 9360 598
rect 9398 201 9404 598
rect 9354 189 9404 201
rect 9520 598 9570 610
rect 9520 201 9526 598
rect 9564 201 9570 598
rect 9520 189 9570 201
rect 9686 598 9736 610
rect 9686 201 9692 598
rect 9730 201 9736 598
rect 9686 189 9736 201
rect 9852 598 9902 610
rect 9852 201 9858 598
rect 9896 201 9902 598
rect 9852 189 9902 201
rect 10018 598 10068 610
rect 10018 201 10024 598
rect 10062 201 10068 598
rect 10018 189 10068 201
rect 10184 598 10234 610
rect 10184 201 10190 598
rect 10228 201 10234 598
rect 10184 189 10234 201
rect 10350 598 10400 610
rect 10350 201 10356 598
rect 10394 201 10400 598
rect 10350 189 10400 201
rect 10516 598 10566 610
rect 10516 201 10522 598
rect 10560 201 10566 598
rect 10516 189 10566 201
rect 10682 598 10732 610
rect 10682 201 10688 598
rect 10726 201 10732 598
rect 10682 189 10732 201
rect 10848 598 10898 610
rect 10848 201 10854 598
rect 10892 201 10898 598
rect 10848 189 10898 201
rect 11014 598 11064 610
rect 11014 201 11020 598
rect 11058 201 11064 598
rect 11014 189 11064 201
rect 11180 598 11230 610
rect 11180 201 11186 598
rect 11224 201 11230 598
rect 11180 189 11230 201
rect 11346 598 11396 610
rect 11346 201 11352 598
rect 11390 201 11396 598
rect 11346 189 11396 201
rect -11396 -201 -11346 -189
rect -11396 -598 -11390 -201
rect -11352 -598 -11346 -201
rect -11396 -610 -11346 -598
rect -11230 -201 -11180 -189
rect -11230 -598 -11224 -201
rect -11186 -598 -11180 -201
rect -11230 -610 -11180 -598
rect -11064 -201 -11014 -189
rect -11064 -598 -11058 -201
rect -11020 -598 -11014 -201
rect -11064 -610 -11014 -598
rect -10898 -201 -10848 -189
rect -10898 -598 -10892 -201
rect -10854 -598 -10848 -201
rect -10898 -610 -10848 -598
rect -10732 -201 -10682 -189
rect -10732 -598 -10726 -201
rect -10688 -598 -10682 -201
rect -10732 -610 -10682 -598
rect -10566 -201 -10516 -189
rect -10566 -598 -10560 -201
rect -10522 -598 -10516 -201
rect -10566 -610 -10516 -598
rect -10400 -201 -10350 -189
rect -10400 -598 -10394 -201
rect -10356 -598 -10350 -201
rect -10400 -610 -10350 -598
rect -10234 -201 -10184 -189
rect -10234 -598 -10228 -201
rect -10190 -598 -10184 -201
rect -10234 -610 -10184 -598
rect -10068 -201 -10018 -189
rect -10068 -598 -10062 -201
rect -10024 -598 -10018 -201
rect -10068 -610 -10018 -598
rect -9902 -201 -9852 -189
rect -9902 -598 -9896 -201
rect -9858 -598 -9852 -201
rect -9902 -610 -9852 -598
rect -9736 -201 -9686 -189
rect -9736 -598 -9730 -201
rect -9692 -598 -9686 -201
rect -9736 -610 -9686 -598
rect -9570 -201 -9520 -189
rect -9570 -598 -9564 -201
rect -9526 -598 -9520 -201
rect -9570 -610 -9520 -598
rect -9404 -201 -9354 -189
rect -9404 -598 -9398 -201
rect -9360 -598 -9354 -201
rect -9404 -610 -9354 -598
rect -9238 -201 -9188 -189
rect -9238 -598 -9232 -201
rect -9194 -598 -9188 -201
rect -9238 -610 -9188 -598
rect -9072 -201 -9022 -189
rect -9072 -598 -9066 -201
rect -9028 -598 -9022 -201
rect -9072 -610 -9022 -598
rect -8906 -201 -8856 -189
rect -8906 -598 -8900 -201
rect -8862 -598 -8856 -201
rect -8906 -610 -8856 -598
rect -8740 -201 -8690 -189
rect -8740 -598 -8734 -201
rect -8696 -598 -8690 -201
rect -8740 -610 -8690 -598
rect -8574 -201 -8524 -189
rect -8574 -598 -8568 -201
rect -8530 -598 -8524 -201
rect -8574 -610 -8524 -598
rect -8408 -201 -8358 -189
rect -8408 -598 -8402 -201
rect -8364 -598 -8358 -201
rect -8408 -610 -8358 -598
rect -8242 -201 -8192 -189
rect -8242 -598 -8236 -201
rect -8198 -598 -8192 -201
rect -8242 -610 -8192 -598
rect -8076 -201 -8026 -189
rect -8076 -598 -8070 -201
rect -8032 -598 -8026 -201
rect -8076 -610 -8026 -598
rect -7910 -201 -7860 -189
rect -7910 -598 -7904 -201
rect -7866 -598 -7860 -201
rect -7910 -610 -7860 -598
rect -7744 -201 -7694 -189
rect -7744 -598 -7738 -201
rect -7700 -598 -7694 -201
rect -7744 -610 -7694 -598
rect -7578 -201 -7528 -189
rect -7578 -598 -7572 -201
rect -7534 -598 -7528 -201
rect -7578 -610 -7528 -598
rect -7412 -201 -7362 -189
rect -7412 -598 -7406 -201
rect -7368 -598 -7362 -201
rect -7412 -610 -7362 -598
rect -7246 -201 -7196 -189
rect -7246 -598 -7240 -201
rect -7202 -598 -7196 -201
rect -7246 -610 -7196 -598
rect -7080 -201 -7030 -189
rect -7080 -598 -7074 -201
rect -7036 -598 -7030 -201
rect -7080 -610 -7030 -598
rect -6914 -201 -6864 -189
rect -6914 -598 -6908 -201
rect -6870 -598 -6864 -201
rect -6914 -610 -6864 -598
rect -6748 -201 -6698 -189
rect -6748 -598 -6742 -201
rect -6704 -598 -6698 -201
rect -6748 -610 -6698 -598
rect -6582 -201 -6532 -189
rect -6582 -598 -6576 -201
rect -6538 -598 -6532 -201
rect -6582 -610 -6532 -598
rect -6416 -201 -6366 -189
rect -6416 -598 -6410 -201
rect -6372 -598 -6366 -201
rect -6416 -610 -6366 -598
rect -6250 -201 -6200 -189
rect -6250 -598 -6244 -201
rect -6206 -598 -6200 -201
rect -6250 -610 -6200 -598
rect -6084 -201 -6034 -189
rect -6084 -598 -6078 -201
rect -6040 -598 -6034 -201
rect -6084 -610 -6034 -598
rect -5918 -201 -5868 -189
rect -5918 -598 -5912 -201
rect -5874 -598 -5868 -201
rect -5918 -610 -5868 -598
rect -5752 -201 -5702 -189
rect -5752 -598 -5746 -201
rect -5708 -598 -5702 -201
rect -5752 -610 -5702 -598
rect -5586 -201 -5536 -189
rect -5586 -598 -5580 -201
rect -5542 -598 -5536 -201
rect -5586 -610 -5536 -598
rect -5420 -201 -5370 -189
rect -5420 -598 -5414 -201
rect -5376 -598 -5370 -201
rect -5420 -610 -5370 -598
rect -5254 -201 -5204 -189
rect -5254 -598 -5248 -201
rect -5210 -598 -5204 -201
rect -5254 -610 -5204 -598
rect -5088 -201 -5038 -189
rect -5088 -598 -5082 -201
rect -5044 -598 -5038 -201
rect -5088 -610 -5038 -598
rect -4922 -201 -4872 -189
rect -4922 -598 -4916 -201
rect -4878 -598 -4872 -201
rect -4922 -610 -4872 -598
rect -4756 -201 -4706 -189
rect -4756 -598 -4750 -201
rect -4712 -598 -4706 -201
rect -4756 -610 -4706 -598
rect -4590 -201 -4540 -189
rect -4590 -598 -4584 -201
rect -4546 -598 -4540 -201
rect -4590 -610 -4540 -598
rect -4424 -201 -4374 -189
rect -4424 -598 -4418 -201
rect -4380 -598 -4374 -201
rect -4424 -610 -4374 -598
rect -4258 -201 -4208 -189
rect -4258 -598 -4252 -201
rect -4214 -598 -4208 -201
rect -4258 -610 -4208 -598
rect -4092 -201 -4042 -189
rect -4092 -598 -4086 -201
rect -4048 -598 -4042 -201
rect -4092 -610 -4042 -598
rect -3926 -201 -3876 -189
rect -3926 -598 -3920 -201
rect -3882 -598 -3876 -201
rect -3926 -610 -3876 -598
rect -3760 -201 -3710 -189
rect -3760 -598 -3754 -201
rect -3716 -598 -3710 -201
rect -3760 -610 -3710 -598
rect -3594 -201 -3544 -189
rect -3594 -598 -3588 -201
rect -3550 -598 -3544 -201
rect -3594 -610 -3544 -598
rect -3428 -201 -3378 -189
rect -3428 -598 -3422 -201
rect -3384 -598 -3378 -201
rect -3428 -610 -3378 -598
rect -3262 -201 -3212 -189
rect -3262 -598 -3256 -201
rect -3218 -598 -3212 -201
rect -3262 -610 -3212 -598
rect -3096 -201 -3046 -189
rect -3096 -598 -3090 -201
rect -3052 -598 -3046 -201
rect -3096 -610 -3046 -598
rect -2930 -201 -2880 -189
rect -2930 -598 -2924 -201
rect -2886 -598 -2880 -201
rect -2930 -610 -2880 -598
rect -2764 -201 -2714 -189
rect -2764 -598 -2758 -201
rect -2720 -598 -2714 -201
rect -2764 -610 -2714 -598
rect -2598 -201 -2548 -189
rect -2598 -598 -2592 -201
rect -2554 -598 -2548 -201
rect -2598 -610 -2548 -598
rect -2432 -201 -2382 -189
rect -2432 -598 -2426 -201
rect -2388 -598 -2382 -201
rect -2432 -610 -2382 -598
rect -2266 -201 -2216 -189
rect -2266 -598 -2260 -201
rect -2222 -598 -2216 -201
rect -2266 -610 -2216 -598
rect -2100 -201 -2050 -189
rect -2100 -598 -2094 -201
rect -2056 -598 -2050 -201
rect -2100 -610 -2050 -598
rect -1934 -201 -1884 -189
rect -1934 -598 -1928 -201
rect -1890 -598 -1884 -201
rect -1934 -610 -1884 -598
rect -1768 -201 -1718 -189
rect -1768 -598 -1762 -201
rect -1724 -598 -1718 -201
rect -1768 -610 -1718 -598
rect -1602 -201 -1552 -189
rect -1602 -598 -1596 -201
rect -1558 -598 -1552 -201
rect -1602 -610 -1552 -598
rect -1436 -201 -1386 -189
rect -1436 -598 -1430 -201
rect -1392 -598 -1386 -201
rect -1436 -610 -1386 -598
rect -1270 -201 -1220 -189
rect -1270 -598 -1264 -201
rect -1226 -598 -1220 -201
rect -1270 -610 -1220 -598
rect -1104 -201 -1054 -189
rect -1104 -598 -1098 -201
rect -1060 -598 -1054 -201
rect -1104 -610 -1054 -598
rect -938 -201 -888 -189
rect -938 -598 -932 -201
rect -894 -598 -888 -201
rect -938 -610 -888 -598
rect -772 -201 -722 -189
rect -772 -598 -766 -201
rect -728 -598 -722 -201
rect -772 -610 -722 -598
rect -606 -201 -556 -189
rect -606 -598 -600 -201
rect -562 -598 -556 -201
rect -606 -610 -556 -598
rect -440 -201 -390 -189
rect -440 -598 -434 -201
rect -396 -598 -390 -201
rect -440 -610 -390 -598
rect -274 -201 -224 -189
rect -274 -598 -268 -201
rect -230 -598 -224 -201
rect -274 -610 -224 -598
rect -108 -201 -58 -189
rect -108 -598 -102 -201
rect -64 -598 -58 -201
rect -108 -610 -58 -598
rect 58 -201 108 -189
rect 58 -598 64 -201
rect 102 -598 108 -201
rect 58 -610 108 -598
rect 224 -201 274 -189
rect 224 -598 230 -201
rect 268 -598 274 -201
rect 224 -610 274 -598
rect 390 -201 440 -189
rect 390 -598 396 -201
rect 434 -598 440 -201
rect 390 -610 440 -598
rect 556 -201 606 -189
rect 556 -598 562 -201
rect 600 -598 606 -201
rect 556 -610 606 -598
rect 722 -201 772 -189
rect 722 -598 728 -201
rect 766 -598 772 -201
rect 722 -610 772 -598
rect 888 -201 938 -189
rect 888 -598 894 -201
rect 932 -598 938 -201
rect 888 -610 938 -598
rect 1054 -201 1104 -189
rect 1054 -598 1060 -201
rect 1098 -598 1104 -201
rect 1054 -610 1104 -598
rect 1220 -201 1270 -189
rect 1220 -598 1226 -201
rect 1264 -598 1270 -201
rect 1220 -610 1270 -598
rect 1386 -201 1436 -189
rect 1386 -598 1392 -201
rect 1430 -598 1436 -201
rect 1386 -610 1436 -598
rect 1552 -201 1602 -189
rect 1552 -598 1558 -201
rect 1596 -598 1602 -201
rect 1552 -610 1602 -598
rect 1718 -201 1768 -189
rect 1718 -598 1724 -201
rect 1762 -598 1768 -201
rect 1718 -610 1768 -598
rect 1884 -201 1934 -189
rect 1884 -598 1890 -201
rect 1928 -598 1934 -201
rect 1884 -610 1934 -598
rect 2050 -201 2100 -189
rect 2050 -598 2056 -201
rect 2094 -598 2100 -201
rect 2050 -610 2100 -598
rect 2216 -201 2266 -189
rect 2216 -598 2222 -201
rect 2260 -598 2266 -201
rect 2216 -610 2266 -598
rect 2382 -201 2432 -189
rect 2382 -598 2388 -201
rect 2426 -598 2432 -201
rect 2382 -610 2432 -598
rect 2548 -201 2598 -189
rect 2548 -598 2554 -201
rect 2592 -598 2598 -201
rect 2548 -610 2598 -598
rect 2714 -201 2764 -189
rect 2714 -598 2720 -201
rect 2758 -598 2764 -201
rect 2714 -610 2764 -598
rect 2880 -201 2930 -189
rect 2880 -598 2886 -201
rect 2924 -598 2930 -201
rect 2880 -610 2930 -598
rect 3046 -201 3096 -189
rect 3046 -598 3052 -201
rect 3090 -598 3096 -201
rect 3046 -610 3096 -598
rect 3212 -201 3262 -189
rect 3212 -598 3218 -201
rect 3256 -598 3262 -201
rect 3212 -610 3262 -598
rect 3378 -201 3428 -189
rect 3378 -598 3384 -201
rect 3422 -598 3428 -201
rect 3378 -610 3428 -598
rect 3544 -201 3594 -189
rect 3544 -598 3550 -201
rect 3588 -598 3594 -201
rect 3544 -610 3594 -598
rect 3710 -201 3760 -189
rect 3710 -598 3716 -201
rect 3754 -598 3760 -201
rect 3710 -610 3760 -598
rect 3876 -201 3926 -189
rect 3876 -598 3882 -201
rect 3920 -598 3926 -201
rect 3876 -610 3926 -598
rect 4042 -201 4092 -189
rect 4042 -598 4048 -201
rect 4086 -598 4092 -201
rect 4042 -610 4092 -598
rect 4208 -201 4258 -189
rect 4208 -598 4214 -201
rect 4252 -598 4258 -201
rect 4208 -610 4258 -598
rect 4374 -201 4424 -189
rect 4374 -598 4380 -201
rect 4418 -598 4424 -201
rect 4374 -610 4424 -598
rect 4540 -201 4590 -189
rect 4540 -598 4546 -201
rect 4584 -598 4590 -201
rect 4540 -610 4590 -598
rect 4706 -201 4756 -189
rect 4706 -598 4712 -201
rect 4750 -598 4756 -201
rect 4706 -610 4756 -598
rect 4872 -201 4922 -189
rect 4872 -598 4878 -201
rect 4916 -598 4922 -201
rect 4872 -610 4922 -598
rect 5038 -201 5088 -189
rect 5038 -598 5044 -201
rect 5082 -598 5088 -201
rect 5038 -610 5088 -598
rect 5204 -201 5254 -189
rect 5204 -598 5210 -201
rect 5248 -598 5254 -201
rect 5204 -610 5254 -598
rect 5370 -201 5420 -189
rect 5370 -598 5376 -201
rect 5414 -598 5420 -201
rect 5370 -610 5420 -598
rect 5536 -201 5586 -189
rect 5536 -598 5542 -201
rect 5580 -598 5586 -201
rect 5536 -610 5586 -598
rect 5702 -201 5752 -189
rect 5702 -598 5708 -201
rect 5746 -598 5752 -201
rect 5702 -610 5752 -598
rect 5868 -201 5918 -189
rect 5868 -598 5874 -201
rect 5912 -598 5918 -201
rect 5868 -610 5918 -598
rect 6034 -201 6084 -189
rect 6034 -598 6040 -201
rect 6078 -598 6084 -201
rect 6034 -610 6084 -598
rect 6200 -201 6250 -189
rect 6200 -598 6206 -201
rect 6244 -598 6250 -201
rect 6200 -610 6250 -598
rect 6366 -201 6416 -189
rect 6366 -598 6372 -201
rect 6410 -598 6416 -201
rect 6366 -610 6416 -598
rect 6532 -201 6582 -189
rect 6532 -598 6538 -201
rect 6576 -598 6582 -201
rect 6532 -610 6582 -598
rect 6698 -201 6748 -189
rect 6698 -598 6704 -201
rect 6742 -598 6748 -201
rect 6698 -610 6748 -598
rect 6864 -201 6914 -189
rect 6864 -598 6870 -201
rect 6908 -598 6914 -201
rect 6864 -610 6914 -598
rect 7030 -201 7080 -189
rect 7030 -598 7036 -201
rect 7074 -598 7080 -201
rect 7030 -610 7080 -598
rect 7196 -201 7246 -189
rect 7196 -598 7202 -201
rect 7240 -598 7246 -201
rect 7196 -610 7246 -598
rect 7362 -201 7412 -189
rect 7362 -598 7368 -201
rect 7406 -598 7412 -201
rect 7362 -610 7412 -598
rect 7528 -201 7578 -189
rect 7528 -598 7534 -201
rect 7572 -598 7578 -201
rect 7528 -610 7578 -598
rect 7694 -201 7744 -189
rect 7694 -598 7700 -201
rect 7738 -598 7744 -201
rect 7694 -610 7744 -598
rect 7860 -201 7910 -189
rect 7860 -598 7866 -201
rect 7904 -598 7910 -201
rect 7860 -610 7910 -598
rect 8026 -201 8076 -189
rect 8026 -598 8032 -201
rect 8070 -598 8076 -201
rect 8026 -610 8076 -598
rect 8192 -201 8242 -189
rect 8192 -598 8198 -201
rect 8236 -598 8242 -201
rect 8192 -610 8242 -598
rect 8358 -201 8408 -189
rect 8358 -598 8364 -201
rect 8402 -598 8408 -201
rect 8358 -610 8408 -598
rect 8524 -201 8574 -189
rect 8524 -598 8530 -201
rect 8568 -598 8574 -201
rect 8524 -610 8574 -598
rect 8690 -201 8740 -189
rect 8690 -598 8696 -201
rect 8734 -598 8740 -201
rect 8690 -610 8740 -598
rect 8856 -201 8906 -189
rect 8856 -598 8862 -201
rect 8900 -598 8906 -201
rect 8856 -610 8906 -598
rect 9022 -201 9072 -189
rect 9022 -598 9028 -201
rect 9066 -598 9072 -201
rect 9022 -610 9072 -598
rect 9188 -201 9238 -189
rect 9188 -598 9194 -201
rect 9232 -598 9238 -201
rect 9188 -610 9238 -598
rect 9354 -201 9404 -189
rect 9354 -598 9360 -201
rect 9398 -598 9404 -201
rect 9354 -610 9404 -598
rect 9520 -201 9570 -189
rect 9520 -598 9526 -201
rect 9564 -598 9570 -201
rect 9520 -610 9570 -598
rect 9686 -201 9736 -189
rect 9686 -598 9692 -201
rect 9730 -598 9736 -201
rect 9686 -610 9736 -598
rect 9852 -201 9902 -189
rect 9852 -598 9858 -201
rect 9896 -598 9902 -201
rect 9852 -610 9902 -598
rect 10018 -201 10068 -189
rect 10018 -598 10024 -201
rect 10062 -598 10068 -201
rect 10018 -610 10068 -598
rect 10184 -201 10234 -189
rect 10184 -598 10190 -201
rect 10228 -598 10234 -201
rect 10184 -610 10234 -598
rect 10350 -201 10400 -189
rect 10350 -598 10356 -201
rect 10394 -598 10400 -201
rect 10350 -610 10400 -598
rect 10516 -201 10566 -189
rect 10516 -598 10522 -201
rect 10560 -598 10566 -201
rect 10516 -610 10566 -598
rect 10682 -201 10732 -189
rect 10682 -598 10688 -201
rect 10726 -598 10732 -201
rect 10682 -610 10732 -598
rect 10848 -201 10898 -189
rect 10848 -598 10854 -201
rect 10892 -598 10898 -201
rect 10848 -610 10898 -598
rect 11014 -201 11064 -189
rect 11014 -598 11020 -201
rect 11058 -598 11064 -201
rect 11014 -610 11064 -598
rect 11180 -201 11230 -189
rect 11180 -598 11186 -201
rect 11224 -598 11230 -201
rect 11180 -610 11230 -598
rect 11346 -201 11396 -189
rect 11346 -598 11352 -201
rect 11390 -598 11396 -201
rect 11346 -610 11396 -598
<< labels >>
rlabel psubdiffcont 0 -729 0 -729 0 B
port 1 nsew
rlabel xpolycontact -11371 581 -11371 581 0 R1_0
port 2 nsew
rlabel xpolycontact -11371 -581 -11371 -581 0 R2_0
port 3 nsew
rlabel xpolycontact -11205 581 -11205 581 0 R1_1
port 4 nsew
rlabel xpolycontact -11205 -581 -11205 -581 0 R2_1
port 5 nsew
rlabel xpolycontact -11039 581 -11039 581 0 R1_2
port 6 nsew
rlabel xpolycontact -11039 -581 -11039 -581 0 R2_2
port 7 nsew
rlabel xpolycontact -10873 581 -10873 581 0 R1_3
port 8 nsew
rlabel xpolycontact -10873 -581 -10873 -581 0 R2_3
port 9 nsew
rlabel xpolycontact -10707 581 -10707 581 0 R1_4
port 10 nsew
rlabel xpolycontact -10707 -581 -10707 -581 0 R2_4
port 11 nsew
rlabel xpolycontact -10541 581 -10541 581 0 R1_5
port 12 nsew
rlabel xpolycontact -10541 -581 -10541 -581 0 R2_5
port 13 nsew
rlabel xpolycontact -10375 581 -10375 581 0 R1_6
port 14 nsew
rlabel xpolycontact -10375 -581 -10375 -581 0 R2_6
port 15 nsew
rlabel xpolycontact -10209 581 -10209 581 0 R1_7
port 16 nsew
rlabel xpolycontact -10209 -581 -10209 -581 0 R2_7
port 17 nsew
rlabel xpolycontact -10043 581 -10043 581 0 R1_8
port 18 nsew
rlabel xpolycontact -10043 -581 -10043 -581 0 R2_8
port 19 nsew
rlabel xpolycontact -9877 581 -9877 581 0 R1_9
port 20 nsew
rlabel xpolycontact -9877 -581 -9877 -581 0 R2_9
port 21 nsew
rlabel xpolycontact -9711 581 -9711 581 0 R1_10
port 22 nsew
rlabel xpolycontact -9711 -581 -9711 -581 0 R2_10
port 23 nsew
rlabel xpolycontact -9545 581 -9545 581 0 R1_11
port 24 nsew
rlabel xpolycontact -9545 -581 -9545 -581 0 R2_11
port 25 nsew
rlabel xpolycontact -9379 581 -9379 581 0 R1_12
port 26 nsew
rlabel xpolycontact -9379 -581 -9379 -581 0 R2_12
port 27 nsew
rlabel xpolycontact -9213 581 -9213 581 0 R1_13
port 28 nsew
rlabel xpolycontact -9213 -581 -9213 -581 0 R2_13
port 29 nsew
rlabel xpolycontact -9047 581 -9047 581 0 R1_14
port 30 nsew
rlabel xpolycontact -9047 -581 -9047 -581 0 R2_14
port 31 nsew
rlabel xpolycontact -8881 581 -8881 581 0 R1_15
port 32 nsew
rlabel xpolycontact -8881 -581 -8881 -581 0 R2_15
port 33 nsew
rlabel xpolycontact -8715 581 -8715 581 0 R1_16
port 34 nsew
rlabel xpolycontact -8715 -581 -8715 -581 0 R2_16
port 35 nsew
rlabel xpolycontact -8549 581 -8549 581 0 R1_17
port 36 nsew
rlabel xpolycontact -8549 -581 -8549 -581 0 R2_17
port 37 nsew
rlabel xpolycontact -8383 581 -8383 581 0 R1_18
port 38 nsew
rlabel xpolycontact -8383 -581 -8383 -581 0 R2_18
port 39 nsew
rlabel xpolycontact -8217 581 -8217 581 0 R1_19
port 40 nsew
rlabel xpolycontact -8217 -581 -8217 -581 0 R2_19
port 41 nsew
rlabel xpolycontact -8051 581 -8051 581 0 R1_20
port 42 nsew
rlabel xpolycontact -8051 -581 -8051 -581 0 R2_20
port 43 nsew
rlabel xpolycontact -7885 581 -7885 581 0 R1_21
port 44 nsew
rlabel xpolycontact -7885 -581 -7885 -581 0 R2_21
port 45 nsew
rlabel xpolycontact -7719 581 -7719 581 0 R1_22
port 46 nsew
rlabel xpolycontact -7719 -581 -7719 -581 0 R2_22
port 47 nsew
rlabel xpolycontact -7553 581 -7553 581 0 R1_23
port 48 nsew
rlabel xpolycontact -7553 -581 -7553 -581 0 R2_23
port 49 nsew
rlabel xpolycontact -7387 581 -7387 581 0 R1_24
port 50 nsew
rlabel xpolycontact -7387 -581 -7387 -581 0 R2_24
port 51 nsew
rlabel xpolycontact -7221 581 -7221 581 0 R1_25
port 52 nsew
rlabel xpolycontact -7221 -581 -7221 -581 0 R2_25
port 53 nsew
rlabel xpolycontact -7055 581 -7055 581 0 R1_26
port 54 nsew
rlabel xpolycontact -7055 -581 -7055 -581 0 R2_26
port 55 nsew
rlabel xpolycontact -6889 581 -6889 581 0 R1_27
port 56 nsew
rlabel xpolycontact -6889 -581 -6889 -581 0 R2_27
port 57 nsew
rlabel xpolycontact -6723 581 -6723 581 0 R1_28
port 58 nsew
rlabel xpolycontact -6723 -581 -6723 -581 0 R2_28
port 59 nsew
rlabel xpolycontact -6557 581 -6557 581 0 R1_29
port 60 nsew
rlabel xpolycontact -6557 -581 -6557 -581 0 R2_29
port 61 nsew
rlabel xpolycontact -6391 581 -6391 581 0 R1_30
port 62 nsew
rlabel xpolycontact -6391 -581 -6391 -581 0 R2_30
port 63 nsew
rlabel xpolycontact -6225 581 -6225 581 0 R1_31
port 64 nsew
rlabel xpolycontact -6225 -581 -6225 -581 0 R2_31
port 65 nsew
rlabel xpolycontact -6059 581 -6059 581 0 R1_32
port 66 nsew
rlabel xpolycontact -6059 -581 -6059 -581 0 R2_32
port 67 nsew
rlabel xpolycontact -5893 581 -5893 581 0 R1_33
port 68 nsew
rlabel xpolycontact -5893 -581 -5893 -581 0 R2_33
port 69 nsew
rlabel xpolycontact -5727 581 -5727 581 0 R1_34
port 70 nsew
rlabel xpolycontact -5727 -581 -5727 -581 0 R2_34
port 71 nsew
rlabel xpolycontact -5561 581 -5561 581 0 R1_35
port 72 nsew
rlabel xpolycontact -5561 -581 -5561 -581 0 R2_35
port 73 nsew
rlabel xpolycontact -5395 581 -5395 581 0 R1_36
port 74 nsew
rlabel xpolycontact -5395 -581 -5395 -581 0 R2_36
port 75 nsew
rlabel xpolycontact -5229 581 -5229 581 0 R1_37
port 76 nsew
rlabel xpolycontact -5229 -581 -5229 -581 0 R2_37
port 77 nsew
rlabel xpolycontact -5063 581 -5063 581 0 R1_38
port 78 nsew
rlabel xpolycontact -5063 -581 -5063 -581 0 R2_38
port 79 nsew
rlabel xpolycontact -4897 581 -4897 581 0 R1_39
port 80 nsew
rlabel xpolycontact -4897 -581 -4897 -581 0 R2_39
port 81 nsew
rlabel xpolycontact -4731 581 -4731 581 0 R1_40
port 82 nsew
rlabel xpolycontact -4731 -581 -4731 -581 0 R2_40
port 83 nsew
rlabel xpolycontact -4565 581 -4565 581 0 R1_41
port 84 nsew
rlabel xpolycontact -4565 -581 -4565 -581 0 R2_41
port 85 nsew
rlabel xpolycontact -4399 581 -4399 581 0 R1_42
port 86 nsew
rlabel xpolycontact -4399 -581 -4399 -581 0 R2_42
port 87 nsew
rlabel xpolycontact -4233 581 -4233 581 0 R1_43
port 88 nsew
rlabel xpolycontact -4233 -581 -4233 -581 0 R2_43
port 89 nsew
rlabel xpolycontact -4067 581 -4067 581 0 R1_44
port 90 nsew
rlabel xpolycontact -4067 -581 -4067 -581 0 R2_44
port 91 nsew
rlabel xpolycontact -3901 581 -3901 581 0 R1_45
port 92 nsew
rlabel xpolycontact -3901 -581 -3901 -581 0 R2_45
port 93 nsew
rlabel xpolycontact -3735 581 -3735 581 0 R1_46
port 94 nsew
rlabel xpolycontact -3735 -581 -3735 -581 0 R2_46
port 95 nsew
rlabel xpolycontact -3569 581 -3569 581 0 R1_47
port 96 nsew
rlabel xpolycontact -3569 -581 -3569 -581 0 R2_47
port 97 nsew
rlabel xpolycontact -3403 581 -3403 581 0 R1_48
port 98 nsew
rlabel xpolycontact -3403 -581 -3403 -581 0 R2_48
port 99 nsew
rlabel xpolycontact -3237 581 -3237 581 0 R1_49
port 100 nsew
rlabel xpolycontact -3237 -581 -3237 -581 0 R2_49
port 101 nsew
rlabel xpolycontact -3071 581 -3071 581 0 R1_50
port 102 nsew
rlabel xpolycontact -3071 -581 -3071 -581 0 R2_50
port 103 nsew
rlabel xpolycontact -2905 581 -2905 581 0 R1_51
port 104 nsew
rlabel xpolycontact -2905 -581 -2905 -581 0 R2_51
port 105 nsew
rlabel xpolycontact -2739 581 -2739 581 0 R1_52
port 106 nsew
rlabel xpolycontact -2739 -581 -2739 -581 0 R2_52
port 107 nsew
rlabel xpolycontact -2573 581 -2573 581 0 R1_53
port 108 nsew
rlabel xpolycontact -2573 -581 -2573 -581 0 R2_53
port 109 nsew
rlabel xpolycontact -2407 581 -2407 581 0 R1_54
port 110 nsew
rlabel xpolycontact -2407 -581 -2407 -581 0 R2_54
port 111 nsew
rlabel xpolycontact -2241 581 -2241 581 0 R1_55
port 112 nsew
rlabel xpolycontact -2241 -581 -2241 -581 0 R2_55
port 113 nsew
rlabel xpolycontact -2075 581 -2075 581 0 R1_56
port 114 nsew
rlabel xpolycontact -2075 -581 -2075 -581 0 R2_56
port 115 nsew
rlabel xpolycontact -1909 581 -1909 581 0 R1_57
port 116 nsew
rlabel xpolycontact -1909 -581 -1909 -581 0 R2_57
port 117 nsew
rlabel xpolycontact -1743 581 -1743 581 0 R1_58
port 118 nsew
rlabel xpolycontact -1743 -581 -1743 -581 0 R2_58
port 119 nsew
rlabel xpolycontact -1577 581 -1577 581 0 R1_59
port 120 nsew
rlabel xpolycontact -1577 -581 -1577 -581 0 R2_59
port 121 nsew
rlabel xpolycontact -1411 581 -1411 581 0 R1_60
port 122 nsew
rlabel xpolycontact -1411 -581 -1411 -581 0 R2_60
port 123 nsew
rlabel xpolycontact -1245 581 -1245 581 0 R1_61
port 124 nsew
rlabel xpolycontact -1245 -581 -1245 -581 0 R2_61
port 125 nsew
rlabel xpolycontact -1079 581 -1079 581 0 R1_62
port 126 nsew
rlabel xpolycontact -1079 -581 -1079 -581 0 R2_62
port 127 nsew
rlabel xpolycontact -913 581 -913 581 0 R1_63
port 128 nsew
rlabel xpolycontact -913 -581 -913 -581 0 R2_63
port 129 nsew
rlabel xpolycontact -747 581 -747 581 0 R1_64
port 130 nsew
rlabel xpolycontact -747 -581 -747 -581 0 R2_64
port 131 nsew
rlabel xpolycontact -581 581 -581 581 0 R1_65
port 132 nsew
rlabel xpolycontact -581 -581 -581 -581 0 R2_65
port 133 nsew
rlabel xpolycontact -415 581 -415 581 0 R1_66
port 134 nsew
rlabel xpolycontact -415 -581 -415 -581 0 R2_66
port 135 nsew
rlabel xpolycontact -249 581 -249 581 0 R1_67
port 136 nsew
rlabel xpolycontact -249 -581 -249 -581 0 R2_67
port 137 nsew
rlabel xpolycontact -83 581 -83 581 0 R1_68
port 138 nsew
rlabel xpolycontact -83 -581 -83 -581 0 R2_68
port 139 nsew
rlabel xpolycontact 83 581 83 581 0 R1_69
port 140 nsew
rlabel xpolycontact 83 -581 83 -581 0 R2_69
port 141 nsew
rlabel xpolycontact 249 581 249 581 0 R1_70
port 142 nsew
rlabel xpolycontact 249 -581 249 -581 0 R2_70
port 143 nsew
rlabel xpolycontact 415 581 415 581 0 R1_71
port 144 nsew
rlabel xpolycontact 415 -581 415 -581 0 R2_71
port 145 nsew
rlabel xpolycontact 581 581 581 581 0 R1_72
port 146 nsew
rlabel xpolycontact 581 -581 581 -581 0 R2_72
port 147 nsew
rlabel xpolycontact 747 581 747 581 0 R1_73
port 148 nsew
rlabel xpolycontact 747 -581 747 -581 0 R2_73
port 149 nsew
rlabel xpolycontact 913 581 913 581 0 R1_74
port 150 nsew
rlabel xpolycontact 913 -581 913 -581 0 R2_74
port 151 nsew
rlabel xpolycontact 1079 581 1079 581 0 R1_75
port 152 nsew
rlabel xpolycontact 1079 -581 1079 -581 0 R2_75
port 153 nsew
rlabel xpolycontact 1245 581 1245 581 0 R1_76
port 154 nsew
rlabel xpolycontact 1245 -581 1245 -581 0 R2_76
port 155 nsew
rlabel xpolycontact 1411 581 1411 581 0 R1_77
port 156 nsew
rlabel xpolycontact 1411 -581 1411 -581 0 R2_77
port 157 nsew
rlabel xpolycontact 1577 581 1577 581 0 R1_78
port 158 nsew
rlabel xpolycontact 1577 -581 1577 -581 0 R2_78
port 159 nsew
rlabel xpolycontact 1743 581 1743 581 0 R1_79
port 160 nsew
rlabel xpolycontact 1743 -581 1743 -581 0 R2_79
port 161 nsew
rlabel xpolycontact 1909 581 1909 581 0 R1_80
port 162 nsew
rlabel xpolycontact 1909 -581 1909 -581 0 R2_80
port 163 nsew
rlabel xpolycontact 2075 581 2075 581 0 R1_81
port 164 nsew
rlabel xpolycontact 2075 -581 2075 -581 0 R2_81
port 165 nsew
rlabel xpolycontact 2241 581 2241 581 0 R1_82
port 166 nsew
rlabel xpolycontact 2241 -581 2241 -581 0 R2_82
port 167 nsew
rlabel xpolycontact 2407 581 2407 581 0 R1_83
port 168 nsew
rlabel xpolycontact 2407 -581 2407 -581 0 R2_83
port 169 nsew
rlabel xpolycontact 2573 581 2573 581 0 R1_84
port 170 nsew
rlabel xpolycontact 2573 -581 2573 -581 0 R2_84
port 171 nsew
rlabel xpolycontact 2739 581 2739 581 0 R1_85
port 172 nsew
rlabel xpolycontact 2739 -581 2739 -581 0 R2_85
port 173 nsew
rlabel xpolycontact 2905 581 2905 581 0 R1_86
port 174 nsew
rlabel xpolycontact 2905 -581 2905 -581 0 R2_86
port 175 nsew
rlabel xpolycontact 3071 581 3071 581 0 R1_87
port 176 nsew
rlabel xpolycontact 3071 -581 3071 -581 0 R2_87
port 177 nsew
rlabel xpolycontact 3237 581 3237 581 0 R1_88
port 178 nsew
rlabel xpolycontact 3237 -581 3237 -581 0 R2_88
port 179 nsew
rlabel xpolycontact 3403 581 3403 581 0 R1_89
port 180 nsew
rlabel xpolycontact 3403 -581 3403 -581 0 R2_89
port 181 nsew
rlabel xpolycontact 3569 581 3569 581 0 R1_90
port 182 nsew
rlabel xpolycontact 3569 -581 3569 -581 0 R2_90
port 183 nsew
rlabel xpolycontact 3735 581 3735 581 0 R1_91
port 184 nsew
rlabel xpolycontact 3735 -581 3735 -581 0 R2_91
port 185 nsew
rlabel xpolycontact 3901 581 3901 581 0 R1_92
port 186 nsew
rlabel xpolycontact 3901 -581 3901 -581 0 R2_92
port 187 nsew
rlabel xpolycontact 4067 581 4067 581 0 R1_93
port 188 nsew
rlabel xpolycontact 4067 -581 4067 -581 0 R2_93
port 189 nsew
rlabel xpolycontact 4233 581 4233 581 0 R1_94
port 190 nsew
rlabel xpolycontact 4233 -581 4233 -581 0 R2_94
port 191 nsew
rlabel xpolycontact 4399 581 4399 581 0 R1_95
port 192 nsew
rlabel xpolycontact 4399 -581 4399 -581 0 R2_95
port 193 nsew
rlabel xpolycontact 4565 581 4565 581 0 R1_96
port 194 nsew
rlabel xpolycontact 4565 -581 4565 -581 0 R2_96
port 195 nsew
rlabel xpolycontact 4731 581 4731 581 0 R1_97
port 196 nsew
rlabel xpolycontact 4731 -581 4731 -581 0 R2_97
port 197 nsew
rlabel xpolycontact 4897 581 4897 581 0 R1_98
port 198 nsew
rlabel xpolycontact 4897 -581 4897 -581 0 R2_98
port 199 nsew
rlabel xpolycontact 5063 581 5063 581 0 R1_99
port 200 nsew
rlabel xpolycontact 5063 -581 5063 -581 0 R2_99
port 201 nsew
rlabel xpolycontact 5229 581 5229 581 0 R1_100
port 202 nsew
rlabel xpolycontact 5229 -581 5229 -581 0 R2_100
port 203 nsew
rlabel xpolycontact 5395 581 5395 581 0 R1_101
port 204 nsew
rlabel xpolycontact 5395 -581 5395 -581 0 R2_101
port 205 nsew
rlabel xpolycontact 5561 581 5561 581 0 R1_102
port 206 nsew
rlabel xpolycontact 5561 -581 5561 -581 0 R2_102
port 207 nsew
rlabel xpolycontact 5727 581 5727 581 0 R1_103
port 208 nsew
rlabel xpolycontact 5727 -581 5727 -581 0 R2_103
port 209 nsew
rlabel xpolycontact 5893 581 5893 581 0 R1_104
port 210 nsew
rlabel xpolycontact 5893 -581 5893 -581 0 R2_104
port 211 nsew
rlabel xpolycontact 6059 581 6059 581 0 R1_105
port 212 nsew
rlabel xpolycontact 6059 -581 6059 -581 0 R2_105
port 213 nsew
rlabel xpolycontact 6225 581 6225 581 0 R1_106
port 214 nsew
rlabel xpolycontact 6225 -581 6225 -581 0 R2_106
port 215 nsew
rlabel xpolycontact 6391 581 6391 581 0 R1_107
port 216 nsew
rlabel xpolycontact 6391 -581 6391 -581 0 R2_107
port 217 nsew
rlabel xpolycontact 6557 581 6557 581 0 R1_108
port 218 nsew
rlabel xpolycontact 6557 -581 6557 -581 0 R2_108
port 219 nsew
rlabel xpolycontact 6723 581 6723 581 0 R1_109
port 220 nsew
rlabel xpolycontact 6723 -581 6723 -581 0 R2_109
port 221 nsew
rlabel xpolycontact 6889 581 6889 581 0 R1_110
port 222 nsew
rlabel xpolycontact 6889 -581 6889 -581 0 R2_110
port 223 nsew
rlabel xpolycontact 7055 581 7055 581 0 R1_111
port 224 nsew
rlabel xpolycontact 7055 -581 7055 -581 0 R2_111
port 225 nsew
rlabel xpolycontact 7221 581 7221 581 0 R1_112
port 226 nsew
rlabel xpolycontact 7221 -581 7221 -581 0 R2_112
port 227 nsew
rlabel xpolycontact 7387 581 7387 581 0 R1_113
port 228 nsew
rlabel xpolycontact 7387 -581 7387 -581 0 R2_113
port 229 nsew
rlabel xpolycontact 7553 581 7553 581 0 R1_114
port 230 nsew
rlabel xpolycontact 7553 -581 7553 -581 0 R2_114
port 231 nsew
rlabel xpolycontact 7719 581 7719 581 0 R1_115
port 232 nsew
rlabel xpolycontact 7719 -581 7719 -581 0 R2_115
port 233 nsew
rlabel xpolycontact 7885 581 7885 581 0 R1_116
port 234 nsew
rlabel xpolycontact 7885 -581 7885 -581 0 R2_116
port 235 nsew
rlabel xpolycontact 8051 581 8051 581 0 R1_117
port 236 nsew
rlabel xpolycontact 8051 -581 8051 -581 0 R2_117
port 237 nsew
rlabel xpolycontact 8217 581 8217 581 0 R1_118
port 238 nsew
rlabel xpolycontact 8217 -581 8217 -581 0 R2_118
port 239 nsew
rlabel xpolycontact 8383 581 8383 581 0 R1_119
port 240 nsew
rlabel xpolycontact 8383 -581 8383 -581 0 R2_119
port 241 nsew
rlabel xpolycontact 8549 581 8549 581 0 R1_120
port 242 nsew
rlabel xpolycontact 8549 -581 8549 -581 0 R2_120
port 243 nsew
rlabel xpolycontact 8715 581 8715 581 0 R1_121
port 244 nsew
rlabel xpolycontact 8715 -581 8715 -581 0 R2_121
port 245 nsew
rlabel xpolycontact 8881 581 8881 581 0 R1_122
port 246 nsew
rlabel xpolycontact 8881 -581 8881 -581 0 R2_122
port 247 nsew
rlabel xpolycontact 9047 581 9047 581 0 R1_123
port 248 nsew
rlabel xpolycontact 9047 -581 9047 -581 0 R2_123
port 249 nsew
rlabel xpolycontact 9213 581 9213 581 0 R1_124
port 250 nsew
rlabel xpolycontact 9213 -581 9213 -581 0 R2_124
port 251 nsew
rlabel xpolycontact 9379 581 9379 581 0 R1_125
port 252 nsew
rlabel xpolycontact 9379 -581 9379 -581 0 R2_125
port 253 nsew
rlabel xpolycontact 9545 581 9545 581 0 R1_126
port 254 nsew
rlabel xpolycontact 9545 -581 9545 -581 0 R2_126
port 255 nsew
rlabel xpolycontact 9711 581 9711 581 0 R1_127
port 256 nsew
rlabel xpolycontact 9711 -581 9711 -581 0 R2_127
port 257 nsew
rlabel xpolycontact 9877 581 9877 581 0 R1_128
port 258 nsew
rlabel xpolycontact 9877 -581 9877 -581 0 R2_128
port 259 nsew
rlabel xpolycontact 10043 581 10043 581 0 R1_129
port 260 nsew
rlabel xpolycontact 10043 -581 10043 -581 0 R2_129
port 261 nsew
rlabel xpolycontact 10209 581 10209 581 0 R1_130
port 262 nsew
rlabel xpolycontact 10209 -581 10209 -581 0 R2_130
port 263 nsew
rlabel xpolycontact 10375 581 10375 581 0 R1_131
port 264 nsew
rlabel xpolycontact 10375 -581 10375 -581 0 R2_131
port 265 nsew
rlabel xpolycontact 10541 581 10541 581 0 R1_132
port 266 nsew
rlabel xpolycontact 10541 -581 10541 -581 0 R2_132
port 267 nsew
rlabel xpolycontact 10707 581 10707 581 0 R1_133
port 268 nsew
rlabel xpolycontact 10707 -581 10707 -581 0 R2_133
port 269 nsew
rlabel xpolycontact 10873 581 10873 581 0 R1_134
port 270 nsew
rlabel xpolycontact 10873 -581 10873 -581 0 R2_134
port 271 nsew
rlabel xpolycontact 11039 581 11039 581 0 R1_135
port 272 nsew
rlabel xpolycontact 11039 -581 11039 -581 0 R2_135
port 273 nsew
rlabel xpolycontact 11205 581 11205 581 0 R1_136
port 274 nsew
rlabel xpolycontact 11205 -581 11205 -581 0 R2_136
port 275 nsew
rlabel xpolycontact 11371 581 11371 581 0 R1_137
port 276 nsew
rlabel xpolycontact 11371 -581 11371 -581 0 R2_137
port 277 nsew
<< properties >>
string FIXED_BBOX -11519 -729 11519 729
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 2 m 1 nx 138 wmin 0.350 lmin 0.50 class resistor rho 2000 val 12.504k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0 doports 1
<< end >>
