magic
tech sky130A
magscale 1 2
timestamp 1757114530
<< metal1 >>
rect 100 8330 365 8735
rect 475 8330 695 8735
rect 810 8330 1030 8735
rect 1140 8330 1360 8735
rect 1475 8330 1695 8735
rect 1805 8330 2025 8735
rect 2140 8330 2360 8735
rect 2470 8330 2690 8735
rect 2800 8330 3020 8735
rect 3135 8330 3355 8735
rect 3465 8330 3685 8735
rect 3800 8330 4020 8735
rect 4130 8330 4350 8735
rect 4460 8330 4680 8735
rect 4795 8330 5015 8735
rect 5125 8330 5345 8735
rect 5460 8330 5680 8735
rect 5790 8330 6010 8735
rect 6125 8330 6345 8735
rect 6455 8330 6675 8735
rect 6785 8330 7005 8735
rect 7120 8330 7340 8735
rect 7450 8330 7670 8735
rect 7780 8330 8000 8735
rect 8115 8330 8335 8735
rect 8445 8330 8665 8735
rect 8780 8330 9000 8735
rect 9110 8330 9330 8735
rect 9440 8330 9660 8735
rect 9770 8330 9990 8735
rect 10105 8330 10325 8735
rect 10440 8330 10660 8735
rect 10770 8330 10990 8735
rect 11100 8330 11320 8735
rect 11435 8330 11655 8735
rect 11765 8330 11985 8735
rect 12095 8330 12315 8735
rect 12430 8330 12650 8735
rect 12760 8330 12980 8735
rect 13095 8330 13315 8735
rect 13425 8330 13645 8735
rect 13760 8330 13980 8735
rect 14090 8330 14310 8735
rect 14420 8330 14640 8735
rect 14755 8330 14975 8735
rect 15085 8330 15305 8735
rect 15420 8330 15640 8735
rect 15750 8330 15970 8735
rect 16080 8330 16300 8735
rect 16415 8330 16635 8735
rect 17080 8330 17300 8735
rect 17410 8330 17630 8735
rect 17740 8330 17960 8735
rect 18075 8330 18295 8735
rect 18405 8330 18625 8735
rect 18740 8330 18960 8735
rect 19070 8330 19290 8735
rect 19400 8330 19620 8735
rect 19735 8330 19955 8735
rect 20065 8330 20285 8735
rect 20400 8330 20620 8735
rect 20730 8330 20950 8735
rect 21060 8330 21280 8735
rect 21395 8330 21615 8735
rect 21725 8330 21945 8735
rect 22060 8330 22280 8735
rect 22390 8330 22610 8735
rect 22720 8330 22940 8735
rect 23055 8330 23315 8735
rect 310 7530 530 7935
rect 640 7530 865 7935
rect 975 7530 1195 7935
rect 1305 7530 1525 7935
rect 1640 7530 1860 7935
rect 1970 7530 2190 7935
rect 2300 7530 2520 7935
rect 2635 7530 2855 7935
rect 2965 7530 3185 7935
rect 3300 7530 3520 7935
rect 3630 7530 3850 7935
rect 3965 7530 4185 7935
rect 4295 7530 4515 7935
rect 4625 7530 4845 7935
rect 4960 7530 5180 7935
rect 5290 7530 5510 7935
rect 5625 7530 5845 7935
rect 5955 7530 6175 7935
rect 6285 7530 6505 7935
rect 6620 7530 6840 7935
rect 6950 7530 7170 7935
rect 7285 7530 7505 7935
rect 7615 7530 7835 7935
rect 7945 7530 8165 7935
rect 8280 7530 8500 7935
rect 8610 7530 8830 7935
rect 8945 7530 9165 7935
rect 9275 7530 9495 7935
rect 9610 7530 9830 7935
rect 9940 7530 10160 7935
rect 10270 7530 10490 7935
rect 10605 7530 10825 7935
rect 10935 7530 11155 7935
rect 11270 7530 11490 7935
rect 11600 7530 11820 7935
rect 11930 7530 12150 7935
rect 12265 7530 12485 7935
rect 12595 7530 12815 7935
rect 12925 7530 13145 7935
rect 13260 7530 13480 7935
rect 13590 7530 13810 7935
rect 13925 7530 14145 7935
rect 14255 7530 14475 7935
rect 14585 7530 14805 7935
rect 14915 7530 15135 7935
rect 15250 7530 15470 7935
rect 15585 7530 15805 7935
rect 15915 7530 16135 7935
rect 16245 7530 16465 7935
rect 16580 7530 16800 7935
rect 16910 7530 17130 7935
rect 17245 7530 17465 7935
rect 17575 7530 17795 7935
rect 17910 7530 18130 7935
rect 18240 7530 18460 7935
rect 18570 7530 18790 7935
rect 18900 7530 19120 7935
rect 19235 7530 19455 7935
rect 19565 7530 19785 7935
rect 19895 7530 20115 7935
rect 20230 7530 20450 7935
rect 20565 7530 20785 7935
rect 20895 7530 21115 7935
rect 21225 7530 21445 7935
rect 21560 7530 21780 7935
rect 21890 7530 22110 7935
rect 22220 7530 22440 7935
rect 22555 7530 22775 7935
rect 22885 7530 23105 7935
use sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4  sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0
timestamp 1757113279
transform 1 0 11707 0 1 8132
box -11572 -782 11572 782
<< end >>
