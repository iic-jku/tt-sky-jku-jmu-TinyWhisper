VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_TinyWhisper
  CLASS BLOCK ;
  FOREIGN tt_um_TinyWhisper ;
  ORIGIN 0.000 0.000 ;
  SIZE 334.880 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 72.000000 ;
    ANTENNADIFFAREA 20.879999 ;
    PORT
      LAYER li1 ;
        RECT 157.565 45.805 157.915 47.965 ;
        RECT 72.835 32.370 73.005 41.410 ;
        RECT 75.415 32.370 75.585 41.410 ;
        RECT 77.995 32.370 78.165 41.410 ;
        RECT 99.485 32.370 99.655 41.410 ;
        RECT 102.065 32.370 102.235 41.410 ;
        RECT 104.645 32.370 104.815 41.410 ;
        RECT 149.150 31.985 150.150 32.155 ;
        RECT 150.440 31.985 151.440 32.155 ;
        RECT 151.730 31.985 152.730 32.155 ;
        RECT 153.020 31.985 154.020 32.155 ;
        RECT 154.310 31.985 155.310 32.155 ;
        RECT 155.600 31.985 156.600 32.155 ;
        RECT 149.150 30.235 150.150 30.405 ;
        RECT 150.440 30.235 151.440 30.405 ;
        RECT 151.730 30.235 152.730 30.405 ;
        RECT 153.020 30.235 154.020 30.405 ;
        RECT 154.310 30.235 155.310 30.405 ;
        RECT 155.600 30.235 156.600 30.405 ;
        RECT 72.835 27.025 73.005 30.065 ;
        RECT 75.415 27.025 75.585 30.065 ;
        RECT 77.995 27.025 78.165 30.065 ;
        RECT 99.485 27.025 99.655 30.065 ;
        RECT 102.065 27.025 102.235 30.065 ;
        RECT 104.645 27.025 104.815 30.065 ;
      LAYER met1 ;
        RECT 157.615 47.900 157.865 47.940 ;
        RECT 157.600 45.875 160.200 47.900 ;
        RECT 157.615 45.835 157.865 45.875 ;
        RECT 72.655 32.370 73.180 41.395 ;
        RECT 75.230 32.370 75.755 41.395 ;
        RECT 77.805 32.370 78.330 41.395 ;
        RECT 99.305 32.370 99.830 41.395 ;
        RECT 101.880 32.370 102.405 41.395 ;
        RECT 104.455 32.370 104.980 41.395 ;
        RECT 149.170 32.145 150.130 32.185 ;
        RECT 150.460 32.145 151.420 32.185 ;
        RECT 151.750 32.145 152.710 32.185 ;
        RECT 153.040 32.145 154.000 32.185 ;
        RECT 154.330 32.145 155.290 32.185 ;
        RECT 155.620 32.145 156.580 32.185 ;
        RECT 149.170 31.955 156.580 32.145 ;
        RECT 149.180 31.470 156.580 31.955 ;
        RECT 146.330 30.920 156.580 31.470 ;
        RECT 149.180 30.435 156.580 30.920 ;
        RECT 149.170 30.245 156.580 30.435 ;
        RECT 149.170 30.205 150.130 30.245 ;
        RECT 150.460 30.205 151.420 30.245 ;
        RECT 151.750 30.205 152.710 30.245 ;
        RECT 153.040 30.205 154.000 30.245 ;
        RECT 154.330 30.205 155.290 30.245 ;
        RECT 155.620 30.205 156.580 30.245 ;
        RECT 72.680 27.045 73.130 30.045 ;
        RECT 75.280 27.045 75.730 30.045 ;
        RECT 77.855 27.045 78.305 30.045 ;
        RECT 99.330 27.045 99.780 30.045 ;
        RECT 101.930 27.045 102.380 30.045 ;
        RECT 104.505 27.045 104.955 30.045 ;
      LAYER met2 ;
        RECT 158.875 45.875 160.200 47.900 ;
        RECT 72.655 32.370 73.180 41.395 ;
        RECT 75.230 32.370 75.755 41.395 ;
        RECT 77.805 32.370 78.330 41.395 ;
        RECT 72.805 31.470 73.030 32.370 ;
        RECT 75.380 31.470 75.605 32.370 ;
        RECT 77.955 31.470 78.180 32.370 ;
        RECT 81.680 31.470 82.105 37.320 ;
        RECT 99.305 32.370 99.830 41.395 ;
        RECT 101.880 32.370 102.405 41.395 ;
        RECT 104.455 32.370 104.980 41.395 ;
        RECT 72.805 30.920 82.105 31.470 ;
        RECT 99.455 31.470 99.680 32.370 ;
        RECT 102.030 31.470 102.255 32.370 ;
        RECT 104.605 31.470 104.830 32.370 ;
        RECT 108.330 31.470 108.755 37.320 ;
        RECT 99.455 30.920 108.755 31.470 ;
        RECT 146.330 30.920 146.880 31.470 ;
        RECT 72.805 30.045 73.030 30.920 ;
        RECT 75.380 30.045 75.605 30.920 ;
        RECT 77.955 30.045 78.180 30.920 ;
        RECT 99.455 30.045 99.680 30.920 ;
        RECT 102.030 30.045 102.255 30.920 ;
        RECT 104.605 30.045 104.830 30.920 ;
        RECT 72.680 27.045 73.130 30.045 ;
        RECT 75.280 27.045 75.730 30.045 ;
        RECT 77.855 27.045 78.305 30.045 ;
        RECT 99.330 27.045 99.780 30.045 ;
        RECT 101.930 27.045 102.380 30.045 ;
        RECT 104.505 27.045 104.955 30.045 ;
      LAYER met3 ;
        RECT 158.875 44.975 174.125 47.900 ;
        RECT 81.675 43.225 174.125 44.975 ;
        RECT 81.680 36.895 82.105 43.225 ;
        RECT 108.330 36.895 108.755 43.225 ;
        RECT 146.280 31.470 146.705 43.225 ;
        RECT 146.280 30.920 146.880 31.470 ;
      LAYER met4 ;
        RECT 168.060 10.740 172.735 47.905 ;
        RECT 149.765 6.065 172.735 10.740 ;
        RECT 149.765 0.390 154.440 6.065 ;
        RECT 151.810 0.000 152.710 0.390 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 72.000000 ;
    ANTENNADIFFAREA 20.879999 ;
    PORT
      LAYER li1 ;
        RECT 86.160 32.370 86.330 41.410 ;
        RECT 88.740 32.370 88.910 41.410 ;
        RECT 91.320 32.370 91.490 41.410 ;
        RECT 112.810 32.370 112.980 41.410 ;
        RECT 115.390 32.370 115.560 41.410 ;
        RECT 117.970 32.370 118.140 41.410 ;
        RECT 162.475 31.985 163.475 32.155 ;
        RECT 163.765 31.985 164.765 32.155 ;
        RECT 165.055 31.985 166.055 32.155 ;
        RECT 166.345 31.985 167.345 32.155 ;
        RECT 167.635 31.985 168.635 32.155 ;
        RECT 168.925 31.985 169.925 32.155 ;
        RECT 162.475 30.235 163.475 30.405 ;
        RECT 163.765 30.235 164.765 30.405 ;
        RECT 165.055 30.235 166.055 30.405 ;
        RECT 166.345 30.235 167.345 30.405 ;
        RECT 167.635 30.235 168.635 30.405 ;
        RECT 168.925 30.235 169.925 30.405 ;
        RECT 86.160 27.025 86.330 30.065 ;
        RECT 88.740 27.025 88.910 30.065 ;
        RECT 91.320 27.025 91.490 30.065 ;
        RECT 112.810 27.025 112.980 30.065 ;
        RECT 115.390 27.025 115.560 30.065 ;
        RECT 117.970 27.025 118.140 30.065 ;
        RECT 157.565 20.580 157.915 22.740 ;
      LAYER met1 ;
        RECT 85.980 32.370 86.505 41.395 ;
        RECT 88.555 32.370 89.080 41.395 ;
        RECT 91.130 32.370 91.655 41.395 ;
        RECT 112.630 32.370 113.155 41.395 ;
        RECT 115.205 32.370 115.730 41.395 ;
        RECT 117.780 32.370 118.305 41.395 ;
        RECT 162.495 32.145 163.455 32.185 ;
        RECT 163.785 32.145 164.745 32.185 ;
        RECT 165.075 32.145 166.035 32.185 ;
        RECT 166.365 32.145 167.325 32.185 ;
        RECT 167.655 32.145 168.615 32.185 ;
        RECT 168.945 32.145 169.905 32.185 ;
        RECT 162.495 31.955 169.905 32.145 ;
        RECT 162.505 31.470 169.905 31.955 ;
        RECT 159.655 30.920 169.905 31.470 ;
        RECT 162.505 30.435 169.905 30.920 ;
        RECT 162.495 30.245 169.905 30.435 ;
        RECT 162.495 30.205 163.455 30.245 ;
        RECT 163.785 30.205 164.745 30.245 ;
        RECT 165.075 30.205 166.035 30.245 ;
        RECT 166.365 30.205 167.325 30.245 ;
        RECT 167.655 30.205 168.615 30.245 ;
        RECT 168.945 30.205 169.905 30.245 ;
        RECT 86.005 27.045 86.455 30.045 ;
        RECT 88.605 27.045 89.055 30.045 ;
        RECT 91.180 27.045 91.630 30.045 ;
        RECT 112.655 27.045 113.105 30.045 ;
        RECT 115.255 27.045 115.705 30.045 ;
        RECT 117.830 27.045 118.280 30.045 ;
        RECT 157.615 22.675 157.865 22.710 ;
        RECT 157.615 20.650 160.200 22.675 ;
        RECT 157.615 20.605 157.865 20.650 ;
      LAYER met2 ;
        RECT 85.980 32.370 86.505 41.395 ;
        RECT 88.555 32.370 89.080 41.395 ;
        RECT 91.130 32.370 91.655 41.395 ;
        RECT 112.630 32.370 113.155 41.395 ;
        RECT 115.205 32.370 115.730 41.395 ;
        RECT 117.780 32.370 118.305 41.395 ;
        RECT 86.130 31.470 86.355 32.370 ;
        RECT 88.705 31.470 88.930 32.370 ;
        RECT 91.280 31.470 91.505 32.370 ;
        RECT 112.780 31.470 113.005 32.370 ;
        RECT 115.355 31.470 115.580 32.370 ;
        RECT 117.930 31.470 118.155 32.370 ;
        RECT 86.130 30.920 95.430 31.470 ;
        RECT 86.130 30.045 86.355 30.920 ;
        RECT 88.705 30.045 88.930 30.920 ;
        RECT 91.280 30.045 91.505 30.920 ;
        RECT 86.005 27.045 86.455 30.045 ;
        RECT 88.605 27.045 89.055 30.045 ;
        RECT 91.180 27.045 91.630 30.045 ;
        RECT 95.005 28.345 95.430 30.920 ;
        RECT 112.780 30.920 122.080 31.470 ;
        RECT 159.655 30.920 160.205 31.470 ;
        RECT 112.780 30.045 113.005 30.920 ;
        RECT 115.355 30.045 115.580 30.920 ;
        RECT 117.930 30.045 118.155 30.920 ;
        RECT 112.655 27.045 113.105 30.045 ;
        RECT 115.255 27.045 115.705 30.045 ;
        RECT 117.830 27.045 118.280 30.045 ;
        RECT 121.655 28.295 122.080 30.920 ;
        RECT 158.875 20.650 160.200 22.675 ;
      LAYER met3 ;
        RECT 159.605 30.920 160.205 31.470 ;
        RECT 95.005 25.250 95.430 28.770 ;
        RECT 121.655 25.250 122.080 28.720 ;
        RECT 159.605 25.250 160.030 30.920 ;
        RECT 95.000 23.575 174.125 25.250 ;
        RECT 158.875 20.650 174.125 23.575 ;
        RECT 164.125 15.825 168.725 20.650 ;
        RECT 130.575 11.225 168.725 15.825 ;
        RECT 130.575 5.870 135.175 11.225 ;
      LAYER met4 ;
        RECT 130.570 5.895 135.180 10.495 ;
        RECT 130.575 0.275 135.175 5.895 ;
        RECT 132.490 0.000 133.390 0.275 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 43.855 45.805 44.205 47.965 ;
      LAYER met1 ;
        RECT 24.240 47.900 26.265 47.930 ;
        RECT 43.905 47.900 44.155 47.940 ;
        RECT 21.070 45.875 44.175 47.900 ;
        RECT 24.240 45.845 26.265 45.875 ;
        RECT 43.905 45.835 44.155 45.875 ;
      LAYER met2 ;
        RECT 21.100 47.900 23.125 47.930 ;
        RECT 12.015 45.875 23.125 47.900 ;
        RECT 12.015 40.445 14.040 45.875 ;
        RECT 21.100 45.845 23.125 45.875 ;
      LAYER met3 ;
        RECT 11.990 40.435 14.065 42.510 ;
        RECT 11.990 27.845 14.065 29.860 ;
      LAYER met4 ;
        RECT 11.985 40.460 14.070 42.485 ;
        RECT 12.015 29.725 14.040 40.460 ;
        RECT 11.990 27.840 14.040 29.725 ;
        RECT 11.990 13.535 14.015 27.840 ;
        RECT 11.990 11.515 114.610 13.535 ;
        RECT 112.590 0.290 114.610 11.515 ;
        RECT 113.170 0.000 114.070 0.290 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 43.855 20.580 44.205 22.740 ;
      LAYER met1 ;
        RECT 43.905 22.675 44.155 22.710 ;
        RECT 21.075 20.650 44.175 22.675 ;
        RECT 32.820 11.215 34.845 20.650 ;
        RECT 43.905 20.605 44.155 20.650 ;
        RECT 32.820 9.190 95.235 11.215 ;
        RECT 93.210 8.675 95.235 9.190 ;
        RECT 93.205 6.580 95.240 8.675 ;
      LAYER met2 ;
        RECT 93.175 6.610 95.270 8.645 ;
        RECT 93.205 6.565 95.240 6.610 ;
      LAYER met3 ;
        RECT 93.180 6.555 95.265 8.640 ;
      LAYER met4 ;
        RECT 93.195 8.615 95.245 8.620 ;
        RECT 93.175 6.580 95.270 8.615 ;
        RECT 93.195 0.125 95.245 6.580 ;
        RECT 93.850 0.000 94.750 0.125 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 48.000000 ;
    PORT
      LAYER li1 ;
        RECT 23.625 31.985 24.625 32.155 ;
        RECT 24.915 31.985 25.915 32.155 ;
        RECT 26.205 31.985 27.205 32.155 ;
        RECT 27.495 31.985 28.495 32.155 ;
        RECT 23.625 30.235 24.625 30.405 ;
        RECT 24.915 30.235 25.915 30.405 ;
        RECT 26.205 30.235 27.205 30.405 ;
        RECT 27.495 30.235 28.495 30.405 ;
      LAYER met1 ;
        RECT 23.645 32.145 24.605 32.185 ;
        RECT 24.935 32.145 25.895 32.185 ;
        RECT 26.225 32.145 27.185 32.185 ;
        RECT 27.515 32.145 28.475 32.185 ;
        RECT 23.645 31.955 28.505 32.145 ;
        RECT 21.100 31.470 21.350 31.475 ;
        RECT 23.655 31.470 28.505 31.955 ;
        RECT 21.100 30.925 28.505 31.470 ;
        RECT 21.105 30.920 28.505 30.925 ;
        RECT 23.655 30.435 28.505 30.920 ;
        RECT 23.645 30.245 28.505 30.435 ;
        RECT 23.645 30.205 24.605 30.245 ;
        RECT 24.935 30.205 25.895 30.245 ;
        RECT 26.225 30.205 27.185 30.245 ;
        RECT 27.515 30.205 28.475 30.245 ;
      LAYER met2 ;
        RECT 21.200 31.470 21.750 31.500 ;
        RECT 16.550 30.920 21.750 31.470 ;
        RECT 16.555 6.520 17.095 30.920 ;
        RECT 21.200 30.890 21.750 30.920 ;
        RECT 16.555 5.980 63.290 6.520 ;
      LAYER met3 ;
        RECT 62.730 6.520 63.270 6.545 ;
        RECT 74.730 6.520 75.270 6.540 ;
        RECT 62.730 5.980 75.270 6.520 ;
        RECT 62.730 5.955 63.270 5.980 ;
        RECT 74.730 5.950 75.270 5.980 ;
      LAYER met4 ;
        RECT 74.725 5.975 75.275 6.515 ;
        RECT 74.730 1.000 75.270 5.975 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 43.025 44.975 158.745 52.795 ;
      LAYER nwell ;
        RECT 21.355 31.295 30.765 42.485 ;
        RECT 32.105 31.295 44.095 42.485 ;
        RECT 45.430 31.295 57.420 42.485 ;
        RECT 58.755 31.295 68.165 42.485 ;
        RECT 69.505 31.295 81.495 42.485 ;
        RECT 82.830 31.295 94.820 42.485 ;
        RECT 96.155 31.295 108.145 42.485 ;
        RECT 109.480 31.295 121.470 42.485 ;
        RECT 122.805 31.295 134.795 42.485 ;
        RECT 136.130 31.295 145.540 42.485 ;
        RECT 146.880 31.295 158.870 42.485 ;
        RECT 160.205 31.295 172.195 42.485 ;
      LAYER pwell ;
        RECT 21.355 25.995 30.765 31.095 ;
        RECT 32.105 25.995 44.095 31.095 ;
        RECT 45.430 25.995 57.420 31.095 ;
        RECT 58.755 25.995 68.165 31.095 ;
        RECT 69.505 25.995 81.495 31.095 ;
        RECT 82.830 25.995 94.820 31.095 ;
        RECT 96.155 25.995 108.145 31.095 ;
        RECT 109.480 25.995 121.470 31.095 ;
        RECT 122.805 25.995 134.795 31.095 ;
        RECT 136.130 25.995 145.540 31.095 ;
        RECT 146.880 25.995 158.870 31.095 ;
        RECT 160.205 25.995 172.195 31.095 ;
        RECT 43.025 15.750 158.745 23.570 ;
      LAYER li1 ;
        RECT 43.205 52.445 158.565 52.615 ;
        RECT 43.205 49.175 43.375 52.445 ;
        RECT 43.855 49.805 44.205 51.965 ;
        RECT 44.685 49.805 45.035 51.965 ;
        RECT 45.515 49.805 45.865 51.965 ;
        RECT 46.345 49.805 46.695 51.965 ;
        RECT 47.175 49.805 47.525 51.965 ;
        RECT 48.005 49.805 48.355 51.965 ;
        RECT 48.835 49.805 49.185 51.965 ;
        RECT 49.665 49.805 50.015 51.965 ;
        RECT 50.495 49.805 50.845 51.965 ;
        RECT 51.325 49.805 51.675 51.965 ;
        RECT 52.155 49.805 52.505 51.965 ;
        RECT 52.985 49.805 53.335 51.965 ;
        RECT 53.815 49.805 54.165 51.965 ;
        RECT 54.645 49.805 54.995 51.965 ;
        RECT 55.475 49.805 55.825 51.965 ;
        RECT 56.305 49.805 56.655 51.965 ;
        RECT 57.135 49.805 57.485 51.965 ;
        RECT 57.965 49.805 58.315 51.965 ;
        RECT 58.795 49.805 59.145 51.965 ;
        RECT 59.625 49.805 59.975 51.965 ;
        RECT 60.455 49.805 60.805 51.965 ;
        RECT 61.285 49.805 61.635 51.965 ;
        RECT 62.115 49.805 62.465 51.965 ;
        RECT 62.945 49.805 63.295 51.965 ;
        RECT 63.775 49.805 64.125 51.965 ;
        RECT 64.605 49.805 64.955 51.965 ;
        RECT 65.435 49.805 65.785 51.965 ;
        RECT 66.265 49.805 66.615 51.965 ;
        RECT 67.095 49.805 67.445 51.965 ;
        RECT 67.925 49.805 68.275 51.965 ;
        RECT 68.755 49.805 69.105 51.965 ;
        RECT 69.585 49.805 69.935 51.965 ;
        RECT 70.415 49.805 70.765 51.965 ;
        RECT 71.245 49.805 71.595 51.965 ;
        RECT 72.075 49.805 72.425 51.965 ;
        RECT 72.905 49.805 73.255 51.965 ;
        RECT 73.735 49.805 74.085 51.965 ;
        RECT 74.565 49.805 74.915 51.965 ;
        RECT 75.395 49.805 75.745 51.965 ;
        RECT 76.225 49.805 76.575 51.965 ;
        RECT 77.055 49.805 77.405 51.965 ;
        RECT 77.885 49.805 78.235 51.965 ;
        RECT 78.715 49.805 79.065 51.965 ;
        RECT 79.545 49.805 79.895 51.965 ;
        RECT 80.375 49.805 80.725 51.965 ;
        RECT 81.205 49.805 81.555 51.965 ;
        RECT 82.035 49.805 82.385 51.965 ;
        RECT 82.865 49.805 83.215 51.965 ;
        RECT 83.695 49.805 84.045 51.965 ;
        RECT 84.525 49.805 84.875 51.965 ;
        RECT 85.355 49.805 85.705 51.965 ;
        RECT 86.185 49.805 86.535 51.965 ;
        RECT 87.015 49.805 87.365 51.965 ;
        RECT 87.845 49.805 88.195 51.965 ;
        RECT 88.675 49.805 89.025 51.965 ;
        RECT 89.505 49.805 89.855 51.965 ;
        RECT 90.335 49.805 90.685 51.965 ;
        RECT 91.165 49.805 91.515 51.965 ;
        RECT 91.995 49.805 92.345 51.965 ;
        RECT 92.825 49.805 93.175 51.965 ;
        RECT 93.655 49.805 94.005 51.965 ;
        RECT 94.485 49.805 94.835 51.965 ;
        RECT 95.315 49.805 95.665 51.965 ;
        RECT 96.145 49.805 96.495 51.965 ;
        RECT 96.975 49.805 97.325 51.965 ;
        RECT 97.805 49.805 98.155 51.965 ;
        RECT 98.635 49.805 98.985 51.965 ;
        RECT 99.465 49.805 99.815 51.965 ;
        RECT 100.295 49.805 100.645 51.965 ;
        RECT 101.125 49.805 101.475 51.965 ;
        RECT 101.955 49.805 102.305 51.965 ;
        RECT 102.785 49.805 103.135 51.965 ;
        RECT 103.615 49.805 103.965 51.965 ;
        RECT 104.445 49.805 104.795 51.965 ;
        RECT 105.275 49.805 105.625 51.965 ;
        RECT 106.105 49.805 106.455 51.965 ;
        RECT 106.935 49.805 107.285 51.965 ;
        RECT 107.765 49.805 108.115 51.965 ;
        RECT 108.595 49.805 108.945 51.965 ;
        RECT 109.425 49.805 109.775 51.965 ;
        RECT 110.255 49.805 110.605 51.965 ;
        RECT 111.085 49.805 111.435 51.965 ;
        RECT 111.915 49.805 112.265 51.965 ;
        RECT 112.745 49.805 113.095 51.965 ;
        RECT 113.575 49.805 113.925 51.965 ;
        RECT 114.405 49.805 114.755 51.965 ;
        RECT 115.235 49.805 115.585 51.965 ;
        RECT 116.065 49.805 116.415 51.965 ;
        RECT 116.895 49.805 117.245 51.965 ;
        RECT 117.725 49.805 118.075 51.965 ;
        RECT 118.555 49.805 118.905 51.965 ;
        RECT 119.385 49.805 119.735 51.965 ;
        RECT 120.215 49.805 120.565 51.965 ;
        RECT 121.045 49.805 121.395 51.965 ;
        RECT 121.875 49.805 122.225 51.965 ;
        RECT 122.705 49.805 123.055 51.965 ;
        RECT 123.535 49.805 123.885 51.965 ;
        RECT 124.365 49.805 124.715 51.965 ;
        RECT 125.195 49.805 125.545 51.965 ;
        RECT 126.025 49.805 126.375 51.965 ;
        RECT 126.855 49.805 127.205 51.965 ;
        RECT 127.685 49.805 128.035 51.965 ;
        RECT 128.515 49.805 128.865 51.965 ;
        RECT 129.345 49.805 129.695 51.965 ;
        RECT 130.175 49.805 130.525 51.965 ;
        RECT 131.005 49.805 131.355 51.965 ;
        RECT 131.835 49.805 132.185 51.965 ;
        RECT 132.665 49.805 133.015 51.965 ;
        RECT 133.495 49.805 133.845 51.965 ;
        RECT 134.325 49.805 134.675 51.965 ;
        RECT 135.155 49.805 135.505 51.965 ;
        RECT 135.985 49.805 136.335 51.965 ;
        RECT 136.815 49.805 137.165 51.965 ;
        RECT 137.645 49.805 137.995 51.965 ;
        RECT 138.475 49.805 138.825 51.965 ;
        RECT 139.305 49.805 139.655 51.965 ;
        RECT 140.135 49.805 140.485 51.965 ;
        RECT 140.965 49.805 141.315 51.965 ;
        RECT 141.795 49.805 142.145 51.965 ;
        RECT 142.625 49.805 142.975 51.965 ;
        RECT 143.455 49.805 143.805 51.965 ;
        RECT 144.285 49.805 144.635 51.965 ;
        RECT 145.115 49.805 145.465 51.965 ;
        RECT 145.945 49.805 146.295 51.965 ;
        RECT 146.775 49.805 147.125 51.965 ;
        RECT 147.605 49.805 147.955 51.965 ;
        RECT 148.435 49.805 148.785 51.965 ;
        RECT 149.265 49.805 149.615 51.965 ;
        RECT 150.095 49.805 150.445 51.965 ;
        RECT 150.925 49.805 151.275 51.965 ;
        RECT 151.755 49.805 152.105 51.965 ;
        RECT 152.585 49.805 152.935 51.965 ;
        RECT 153.415 49.805 153.765 51.965 ;
        RECT 154.245 49.805 154.595 51.965 ;
        RECT 155.075 49.805 155.425 51.965 ;
        RECT 155.905 49.805 156.255 51.965 ;
        RECT 156.735 49.805 157.085 51.965 ;
        RECT 157.565 49.805 157.915 51.965 ;
        RECT 43.025 48.550 43.550 49.175 ;
        RECT 43.205 45.325 43.375 48.550 ;
        RECT 44.685 45.805 45.035 47.965 ;
        RECT 45.515 45.805 45.865 47.965 ;
        RECT 46.345 45.805 46.695 47.965 ;
        RECT 47.175 45.805 47.525 47.965 ;
        RECT 48.005 45.805 48.355 47.965 ;
        RECT 48.835 45.805 49.185 47.965 ;
        RECT 49.665 45.805 50.015 47.965 ;
        RECT 50.495 45.805 50.845 47.965 ;
        RECT 51.325 45.805 51.675 47.965 ;
        RECT 52.155 45.805 52.505 47.965 ;
        RECT 52.985 45.805 53.335 47.965 ;
        RECT 53.815 45.805 54.165 47.965 ;
        RECT 54.645 45.805 54.995 47.965 ;
        RECT 55.475 45.805 55.825 47.965 ;
        RECT 56.305 45.805 56.655 47.965 ;
        RECT 57.135 45.805 57.485 47.965 ;
        RECT 57.965 45.805 58.315 47.965 ;
        RECT 58.795 45.805 59.145 47.965 ;
        RECT 59.625 45.805 59.975 47.965 ;
        RECT 60.455 45.805 60.805 47.965 ;
        RECT 61.285 45.805 61.635 47.965 ;
        RECT 62.115 45.805 62.465 47.965 ;
        RECT 62.945 45.805 63.295 47.965 ;
        RECT 63.775 45.805 64.125 47.965 ;
        RECT 64.605 45.805 64.955 47.965 ;
        RECT 65.435 45.805 65.785 47.965 ;
        RECT 66.265 45.805 66.615 47.965 ;
        RECT 67.095 45.805 67.445 47.965 ;
        RECT 67.925 45.805 68.275 47.965 ;
        RECT 68.755 45.805 69.105 47.965 ;
        RECT 69.585 45.805 69.935 47.965 ;
        RECT 70.415 45.805 70.765 47.965 ;
        RECT 71.245 45.805 71.595 47.965 ;
        RECT 72.075 45.805 72.425 47.965 ;
        RECT 72.905 45.805 73.255 47.965 ;
        RECT 73.735 45.805 74.085 47.965 ;
        RECT 74.565 45.805 74.915 47.965 ;
        RECT 75.395 45.805 75.745 47.965 ;
        RECT 76.225 45.805 76.575 47.965 ;
        RECT 77.055 45.805 77.405 47.965 ;
        RECT 77.885 45.805 78.235 47.965 ;
        RECT 78.715 45.805 79.065 47.965 ;
        RECT 79.545 45.805 79.895 47.965 ;
        RECT 80.375 45.805 80.725 47.965 ;
        RECT 81.205 45.805 81.555 47.965 ;
        RECT 82.035 45.805 82.385 47.965 ;
        RECT 82.865 45.805 83.215 47.965 ;
        RECT 83.695 45.805 84.045 47.965 ;
        RECT 84.525 45.805 84.875 47.965 ;
        RECT 85.355 45.805 85.705 47.965 ;
        RECT 86.185 45.805 86.535 47.965 ;
        RECT 87.015 45.805 87.365 47.965 ;
        RECT 87.845 45.805 88.195 47.965 ;
        RECT 88.675 45.805 89.025 47.965 ;
        RECT 89.505 45.805 89.855 47.965 ;
        RECT 90.335 45.805 90.685 47.965 ;
        RECT 91.165 45.805 91.515 47.965 ;
        RECT 91.995 45.805 92.345 47.965 ;
        RECT 92.825 45.805 93.175 47.965 ;
        RECT 93.655 45.805 94.005 47.965 ;
        RECT 94.485 45.805 94.835 47.965 ;
        RECT 95.315 45.805 95.665 47.965 ;
        RECT 96.145 45.805 96.495 47.965 ;
        RECT 96.975 45.805 97.325 47.965 ;
        RECT 97.805 45.805 98.155 47.965 ;
        RECT 98.635 45.805 98.985 47.965 ;
        RECT 99.465 45.805 99.815 47.965 ;
        RECT 100.295 45.805 100.645 47.965 ;
        RECT 101.125 45.805 101.475 47.965 ;
        RECT 101.955 45.805 102.305 47.965 ;
        RECT 102.785 45.805 103.135 47.965 ;
        RECT 103.615 45.805 103.965 47.965 ;
        RECT 104.445 45.805 104.795 47.965 ;
        RECT 105.275 45.805 105.625 47.965 ;
        RECT 106.105 45.805 106.455 47.965 ;
        RECT 106.935 45.805 107.285 47.965 ;
        RECT 107.765 45.805 108.115 47.965 ;
        RECT 108.595 45.805 108.945 47.965 ;
        RECT 109.425 45.805 109.775 47.965 ;
        RECT 110.255 45.805 110.605 47.965 ;
        RECT 111.085 45.805 111.435 47.965 ;
        RECT 111.915 45.805 112.265 47.965 ;
        RECT 112.745 45.805 113.095 47.965 ;
        RECT 113.575 45.805 113.925 47.965 ;
        RECT 114.405 45.805 114.755 47.965 ;
        RECT 115.235 45.805 115.585 47.965 ;
        RECT 116.065 45.805 116.415 47.965 ;
        RECT 116.895 45.805 117.245 47.965 ;
        RECT 117.725 45.805 118.075 47.965 ;
        RECT 118.555 45.805 118.905 47.965 ;
        RECT 119.385 45.805 119.735 47.965 ;
        RECT 120.215 45.805 120.565 47.965 ;
        RECT 121.045 45.805 121.395 47.965 ;
        RECT 121.875 45.805 122.225 47.965 ;
        RECT 122.705 45.805 123.055 47.965 ;
        RECT 123.535 45.805 123.885 47.965 ;
        RECT 124.365 45.805 124.715 47.965 ;
        RECT 125.195 45.805 125.545 47.965 ;
        RECT 126.025 45.805 126.375 47.965 ;
        RECT 126.855 45.805 127.205 47.965 ;
        RECT 127.685 45.805 128.035 47.965 ;
        RECT 128.515 45.805 128.865 47.965 ;
        RECT 129.345 45.805 129.695 47.965 ;
        RECT 130.175 45.805 130.525 47.965 ;
        RECT 131.005 45.805 131.355 47.965 ;
        RECT 131.835 45.805 132.185 47.965 ;
        RECT 132.665 45.805 133.015 47.965 ;
        RECT 133.495 45.805 133.845 47.965 ;
        RECT 134.325 45.805 134.675 47.965 ;
        RECT 135.155 45.805 135.505 47.965 ;
        RECT 135.985 45.805 136.335 47.965 ;
        RECT 136.815 45.805 137.165 47.965 ;
        RECT 137.645 45.805 137.995 47.965 ;
        RECT 138.475 45.805 138.825 47.965 ;
        RECT 139.305 45.805 139.655 47.965 ;
        RECT 140.135 45.805 140.485 47.965 ;
        RECT 140.965 45.805 141.315 47.965 ;
        RECT 141.795 45.805 142.145 47.965 ;
        RECT 142.625 45.805 142.975 47.965 ;
        RECT 143.455 45.805 143.805 47.965 ;
        RECT 144.285 45.805 144.635 47.965 ;
        RECT 145.115 45.805 145.465 47.965 ;
        RECT 145.945 45.805 146.295 47.965 ;
        RECT 146.775 45.805 147.125 47.965 ;
        RECT 147.605 45.805 147.955 47.965 ;
        RECT 148.435 45.805 148.785 47.965 ;
        RECT 149.265 45.805 149.615 47.965 ;
        RECT 150.095 45.805 150.445 47.965 ;
        RECT 150.925 45.805 151.275 47.965 ;
        RECT 151.755 45.805 152.105 47.965 ;
        RECT 152.585 45.805 152.935 47.965 ;
        RECT 153.415 45.805 153.765 47.965 ;
        RECT 154.245 45.805 154.595 47.965 ;
        RECT 155.075 45.805 155.425 47.965 ;
        RECT 155.905 45.805 156.255 47.965 ;
        RECT 156.735 45.805 157.085 47.965 ;
        RECT 158.395 45.325 158.565 52.445 ;
        RECT 43.205 45.155 158.565 45.325 ;
        RECT 21.535 42.135 30.585 42.305 ;
        RECT 21.535 41.320 21.705 42.135 ;
        RECT 22.335 41.625 23.335 41.795 ;
        RECT 28.785 41.625 29.785 41.795 ;
        RECT 21.505 32.445 21.705 41.320 ;
        RECT 21.535 31.645 21.705 32.445 ;
        RECT 22.105 32.370 22.275 41.410 ;
        RECT 23.395 32.370 23.565 41.410 ;
        RECT 24.685 32.370 24.855 41.410 ;
        RECT 25.975 32.370 26.145 41.410 ;
        RECT 27.265 32.370 27.435 41.410 ;
        RECT 28.555 32.370 28.725 41.410 ;
        RECT 29.845 32.370 30.015 41.410 ;
        RECT 30.415 41.320 30.585 42.135 ;
        RECT 32.285 42.135 43.915 42.305 ;
        RECT 32.285 41.320 32.455 42.135 ;
        RECT 33.085 41.625 34.085 41.795 ;
        RECT 42.115 41.625 43.115 41.795 ;
        RECT 30.405 32.445 30.605 41.320 ;
        RECT 32.255 32.445 32.455 41.320 ;
        RECT 30.415 31.645 30.585 32.445 ;
        RECT 21.535 31.475 30.585 31.645 ;
        RECT 32.285 31.645 32.455 32.445 ;
        RECT 32.855 32.370 33.025 41.410 ;
        RECT 34.145 32.370 34.315 41.410 ;
        RECT 35.435 32.370 35.605 41.410 ;
        RECT 36.725 32.370 36.895 41.410 ;
        RECT 38.015 32.370 38.185 41.410 ;
        RECT 39.305 32.370 39.475 41.410 ;
        RECT 40.595 32.370 40.765 41.410 ;
        RECT 41.885 32.370 42.055 41.410 ;
        RECT 43.175 32.370 43.345 41.410 ;
        RECT 43.745 41.320 43.915 42.135 ;
        RECT 45.610 42.135 57.240 42.305 ;
        RECT 45.610 41.320 45.780 42.135 ;
        RECT 46.410 41.625 47.410 41.795 ;
        RECT 55.440 41.625 56.440 41.795 ;
        RECT 43.730 32.445 43.930 41.320 ;
        RECT 45.580 32.445 45.780 41.320 ;
        RECT 34.375 31.985 35.375 32.155 ;
        RECT 35.665 31.985 36.665 32.155 ;
        RECT 36.955 31.985 37.955 32.155 ;
        RECT 38.245 31.985 39.245 32.155 ;
        RECT 39.535 31.985 40.535 32.155 ;
        RECT 40.825 31.985 41.825 32.155 ;
        RECT 43.745 31.645 43.915 32.445 ;
        RECT 32.285 31.475 43.915 31.645 ;
        RECT 45.610 31.645 45.780 32.445 ;
        RECT 46.180 32.370 46.350 41.410 ;
        RECT 47.470 32.370 47.640 41.410 ;
        RECT 48.760 32.370 48.930 41.410 ;
        RECT 50.050 32.370 50.220 41.410 ;
        RECT 51.340 32.370 51.510 41.410 ;
        RECT 52.630 32.370 52.800 41.410 ;
        RECT 53.920 32.370 54.090 41.410 ;
        RECT 55.210 32.370 55.380 41.410 ;
        RECT 56.500 32.370 56.670 41.410 ;
        RECT 57.070 41.320 57.240 42.135 ;
        RECT 58.935 42.135 67.985 42.305 ;
        RECT 58.935 41.320 59.105 42.135 ;
        RECT 59.735 41.625 60.735 41.795 ;
        RECT 66.185 41.625 67.185 41.795 ;
        RECT 57.055 32.445 57.255 41.320 ;
        RECT 58.905 32.445 59.105 41.320 ;
        RECT 47.700 31.985 48.700 32.155 ;
        RECT 48.990 31.985 49.990 32.155 ;
        RECT 50.280 31.985 51.280 32.155 ;
        RECT 51.570 31.985 52.570 32.155 ;
        RECT 52.860 31.985 53.860 32.155 ;
        RECT 54.150 31.985 55.150 32.155 ;
        RECT 57.070 31.645 57.240 32.445 ;
        RECT 45.610 31.475 57.240 31.645 ;
        RECT 58.935 31.645 59.105 32.445 ;
        RECT 59.505 32.370 59.675 41.410 ;
        RECT 60.795 32.370 60.965 41.410 ;
        RECT 62.085 32.370 62.255 41.410 ;
        RECT 63.375 32.370 63.545 41.410 ;
        RECT 64.665 32.370 64.835 41.410 ;
        RECT 65.955 32.370 66.125 41.410 ;
        RECT 67.245 32.370 67.415 41.410 ;
        RECT 67.815 41.320 67.985 42.135 ;
        RECT 69.685 42.135 81.315 42.305 ;
        RECT 69.685 41.320 69.855 42.135 ;
        RECT 70.485 41.625 71.485 41.795 ;
        RECT 79.515 41.625 80.515 41.795 ;
        RECT 67.805 32.445 68.005 41.320 ;
        RECT 69.655 32.445 69.855 41.320 ;
        RECT 61.025 31.985 62.025 32.155 ;
        RECT 62.315 31.985 63.315 32.155 ;
        RECT 63.605 31.985 64.605 32.155 ;
        RECT 64.895 31.985 65.895 32.155 ;
        RECT 67.815 31.645 67.985 32.445 ;
        RECT 58.935 31.475 67.985 31.645 ;
        RECT 69.685 31.645 69.855 32.445 ;
        RECT 70.255 32.370 70.425 41.410 ;
        RECT 71.545 32.370 71.715 41.410 ;
        RECT 74.125 32.370 74.295 41.410 ;
        RECT 76.705 32.370 76.875 41.410 ;
        RECT 79.285 32.370 79.455 41.410 ;
        RECT 80.575 32.370 80.745 41.410 ;
        RECT 81.145 41.320 81.315 42.135 ;
        RECT 83.010 42.135 94.640 42.305 ;
        RECT 83.010 41.320 83.180 42.135 ;
        RECT 83.810 41.625 84.810 41.795 ;
        RECT 92.840 41.625 93.840 41.795 ;
        RECT 81.130 32.445 81.330 41.320 ;
        RECT 82.980 32.445 83.180 41.320 ;
        RECT 71.775 31.985 72.775 32.155 ;
        RECT 73.065 31.985 74.065 32.155 ;
        RECT 74.355 31.985 75.355 32.155 ;
        RECT 75.645 31.985 76.645 32.155 ;
        RECT 76.935 31.985 77.935 32.155 ;
        RECT 78.225 31.985 79.225 32.155 ;
        RECT 81.145 31.645 81.315 32.445 ;
        RECT 69.685 31.475 81.315 31.645 ;
        RECT 83.010 31.645 83.180 32.445 ;
        RECT 83.580 32.370 83.750 41.410 ;
        RECT 84.870 32.370 85.040 41.410 ;
        RECT 87.450 32.370 87.620 41.410 ;
        RECT 90.030 32.370 90.200 41.410 ;
        RECT 92.610 32.370 92.780 41.410 ;
        RECT 93.900 32.370 94.070 41.410 ;
        RECT 94.470 41.320 94.640 42.135 ;
        RECT 96.335 42.135 107.965 42.305 ;
        RECT 96.335 41.320 96.505 42.135 ;
        RECT 97.135 41.625 98.135 41.795 ;
        RECT 106.165 41.625 107.165 41.795 ;
        RECT 94.455 32.445 94.655 41.320 ;
        RECT 96.305 32.445 96.505 41.320 ;
        RECT 85.100 31.985 86.100 32.155 ;
        RECT 86.390 31.985 87.390 32.155 ;
        RECT 87.680 31.985 88.680 32.155 ;
        RECT 88.970 31.985 89.970 32.155 ;
        RECT 90.260 31.985 91.260 32.155 ;
        RECT 91.550 31.985 92.550 32.155 ;
        RECT 94.470 31.645 94.640 32.445 ;
        RECT 83.010 31.475 94.640 31.645 ;
        RECT 96.335 31.645 96.505 32.445 ;
        RECT 96.905 32.370 97.075 41.410 ;
        RECT 98.195 32.370 98.365 41.410 ;
        RECT 100.775 32.370 100.945 41.410 ;
        RECT 103.355 32.370 103.525 41.410 ;
        RECT 105.935 32.370 106.105 41.410 ;
        RECT 107.225 32.370 107.395 41.410 ;
        RECT 107.795 41.320 107.965 42.135 ;
        RECT 109.660 42.135 121.290 42.305 ;
        RECT 109.660 41.320 109.830 42.135 ;
        RECT 110.460 41.625 111.460 41.795 ;
        RECT 119.490 41.625 120.490 41.795 ;
        RECT 107.780 32.445 107.980 41.320 ;
        RECT 109.630 32.445 109.830 41.320 ;
        RECT 98.425 31.985 99.425 32.155 ;
        RECT 99.715 31.985 100.715 32.155 ;
        RECT 101.005 31.985 102.005 32.155 ;
        RECT 102.295 31.985 103.295 32.155 ;
        RECT 103.585 31.985 104.585 32.155 ;
        RECT 104.875 31.985 105.875 32.155 ;
        RECT 107.795 31.645 107.965 32.445 ;
        RECT 96.335 31.475 107.965 31.645 ;
        RECT 109.660 31.645 109.830 32.445 ;
        RECT 110.230 32.370 110.400 41.410 ;
        RECT 111.520 32.370 111.690 41.410 ;
        RECT 114.100 32.370 114.270 41.410 ;
        RECT 116.680 32.370 116.850 41.410 ;
        RECT 119.260 32.370 119.430 41.410 ;
        RECT 120.550 32.370 120.720 41.410 ;
        RECT 121.120 41.320 121.290 42.135 ;
        RECT 122.985 42.135 134.615 42.305 ;
        RECT 122.985 41.320 123.155 42.135 ;
        RECT 123.785 41.625 124.785 41.795 ;
        RECT 132.815 41.625 133.815 41.795 ;
        RECT 121.105 32.445 121.305 41.320 ;
        RECT 122.955 32.445 123.155 41.320 ;
        RECT 111.750 31.985 112.750 32.155 ;
        RECT 113.040 31.985 114.040 32.155 ;
        RECT 114.330 31.985 115.330 32.155 ;
        RECT 115.620 31.985 116.620 32.155 ;
        RECT 116.910 31.985 117.910 32.155 ;
        RECT 118.200 31.985 119.200 32.155 ;
        RECT 121.120 31.645 121.290 32.445 ;
        RECT 109.660 31.475 121.290 31.645 ;
        RECT 122.985 31.645 123.155 32.445 ;
        RECT 123.555 32.370 123.725 41.410 ;
        RECT 124.845 32.370 125.015 41.410 ;
        RECT 126.135 32.370 126.305 41.410 ;
        RECT 127.425 32.370 127.595 41.410 ;
        RECT 128.715 32.370 128.885 41.410 ;
        RECT 130.005 32.370 130.175 41.410 ;
        RECT 131.295 32.370 131.465 41.410 ;
        RECT 132.585 32.370 132.755 41.410 ;
        RECT 133.875 32.370 134.045 41.410 ;
        RECT 134.445 41.320 134.615 42.135 ;
        RECT 136.310 42.135 145.360 42.305 ;
        RECT 136.310 41.320 136.480 42.135 ;
        RECT 137.110 41.625 138.110 41.795 ;
        RECT 143.560 41.625 144.560 41.795 ;
        RECT 134.430 32.445 134.630 41.320 ;
        RECT 136.280 32.445 136.480 41.320 ;
        RECT 125.075 31.985 126.075 32.155 ;
        RECT 126.365 31.985 127.365 32.155 ;
        RECT 127.655 31.985 128.655 32.155 ;
        RECT 128.945 31.985 129.945 32.155 ;
        RECT 130.235 31.985 131.235 32.155 ;
        RECT 131.525 31.985 132.525 32.155 ;
        RECT 134.445 31.645 134.615 32.445 ;
        RECT 122.985 31.475 134.615 31.645 ;
        RECT 136.310 31.645 136.480 32.445 ;
        RECT 136.880 32.370 137.050 41.410 ;
        RECT 138.170 32.370 138.340 41.410 ;
        RECT 139.460 32.370 139.630 41.410 ;
        RECT 140.750 32.370 140.920 41.410 ;
        RECT 142.040 32.370 142.210 41.410 ;
        RECT 143.330 32.370 143.500 41.410 ;
        RECT 144.620 32.370 144.790 41.410 ;
        RECT 145.190 41.320 145.360 42.135 ;
        RECT 147.060 42.135 158.690 42.305 ;
        RECT 147.060 41.320 147.230 42.135 ;
        RECT 147.860 41.625 148.860 41.795 ;
        RECT 156.890 41.625 157.890 41.795 ;
        RECT 145.180 32.445 145.380 41.320 ;
        RECT 147.030 32.445 147.230 41.320 ;
        RECT 138.400 31.985 139.400 32.155 ;
        RECT 139.690 31.985 140.690 32.155 ;
        RECT 140.980 31.985 141.980 32.155 ;
        RECT 142.270 31.985 143.270 32.155 ;
        RECT 145.190 31.645 145.360 32.445 ;
        RECT 136.310 31.475 145.360 31.645 ;
        RECT 147.060 31.645 147.230 32.445 ;
        RECT 147.630 32.370 147.800 41.410 ;
        RECT 148.920 32.370 149.090 41.410 ;
        RECT 150.210 32.370 150.380 41.410 ;
        RECT 151.500 32.370 151.670 41.410 ;
        RECT 152.790 32.370 152.960 41.410 ;
        RECT 154.080 32.370 154.250 41.410 ;
        RECT 155.370 32.370 155.540 41.410 ;
        RECT 156.660 32.370 156.830 41.410 ;
        RECT 157.950 32.370 158.120 41.410 ;
        RECT 158.520 41.320 158.690 42.135 ;
        RECT 160.385 42.135 172.015 42.305 ;
        RECT 160.385 41.320 160.555 42.135 ;
        RECT 161.185 41.625 162.185 41.795 ;
        RECT 170.215 41.625 171.215 41.795 ;
        RECT 158.505 32.445 158.705 41.320 ;
        RECT 160.355 32.445 160.555 41.320 ;
        RECT 158.520 31.645 158.690 32.445 ;
        RECT 147.060 31.475 158.690 31.645 ;
        RECT 160.385 31.645 160.555 32.445 ;
        RECT 160.955 32.370 161.125 41.410 ;
        RECT 162.245 32.370 162.415 41.410 ;
        RECT 163.535 32.370 163.705 41.410 ;
        RECT 164.825 32.370 164.995 41.410 ;
        RECT 166.115 32.370 166.285 41.410 ;
        RECT 167.405 32.370 167.575 41.410 ;
        RECT 168.695 32.370 168.865 41.410 ;
        RECT 169.985 32.370 170.155 41.410 ;
        RECT 171.275 32.370 171.445 41.410 ;
        RECT 171.845 41.320 172.015 42.135 ;
        RECT 171.830 32.445 172.030 41.320 ;
        RECT 171.845 31.645 172.015 32.445 ;
        RECT 160.385 31.475 172.015 31.645 ;
        RECT 21.535 30.745 30.585 30.915 ;
        RECT 21.535 29.995 21.705 30.745 ;
        RECT 21.505 27.095 21.705 29.995 ;
        RECT 21.535 26.345 21.705 27.095 ;
        RECT 22.105 27.025 22.275 30.065 ;
        RECT 23.395 27.025 23.565 30.065 ;
        RECT 24.685 27.025 24.855 30.065 ;
        RECT 25.975 27.025 26.145 30.065 ;
        RECT 27.265 27.025 27.435 30.065 ;
        RECT 28.555 27.025 28.725 30.065 ;
        RECT 29.845 27.025 30.015 30.065 ;
        RECT 30.415 29.995 30.585 30.745 ;
        RECT 32.285 30.745 43.915 30.915 ;
        RECT 32.285 29.995 32.455 30.745 ;
        RECT 34.375 30.235 35.375 30.405 ;
        RECT 35.665 30.235 36.665 30.405 ;
        RECT 36.955 30.235 37.955 30.405 ;
        RECT 38.245 30.235 39.245 30.405 ;
        RECT 39.535 30.235 40.535 30.405 ;
        RECT 40.825 30.235 41.825 30.405 ;
        RECT 30.405 27.095 30.605 29.995 ;
        RECT 32.255 27.095 32.455 29.995 ;
        RECT 22.335 26.685 23.335 26.855 ;
        RECT 28.785 26.685 29.785 26.855 ;
        RECT 30.415 26.345 30.585 27.095 ;
        RECT 21.535 26.175 30.585 26.345 ;
        RECT 32.285 26.345 32.455 27.095 ;
        RECT 32.855 27.025 33.025 30.065 ;
        RECT 34.145 27.025 34.315 30.065 ;
        RECT 35.435 27.025 35.605 30.065 ;
        RECT 36.725 27.025 36.895 30.065 ;
        RECT 38.015 27.025 38.185 30.065 ;
        RECT 39.305 27.025 39.475 30.065 ;
        RECT 40.595 27.025 40.765 30.065 ;
        RECT 41.885 27.025 42.055 30.065 ;
        RECT 43.175 27.025 43.345 30.065 ;
        RECT 43.745 29.995 43.915 30.745 ;
        RECT 45.610 30.745 57.240 30.915 ;
        RECT 45.610 29.995 45.780 30.745 ;
        RECT 47.700 30.235 48.700 30.405 ;
        RECT 48.990 30.235 49.990 30.405 ;
        RECT 50.280 30.235 51.280 30.405 ;
        RECT 51.570 30.235 52.570 30.405 ;
        RECT 52.860 30.235 53.860 30.405 ;
        RECT 54.150 30.235 55.150 30.405 ;
        RECT 43.730 27.095 43.930 29.995 ;
        RECT 45.580 27.095 45.780 29.995 ;
        RECT 33.085 26.685 34.085 26.855 ;
        RECT 42.115 26.685 43.115 26.855 ;
        RECT 43.745 26.345 43.915 27.095 ;
        RECT 32.285 26.175 43.915 26.345 ;
        RECT 45.610 26.345 45.780 27.095 ;
        RECT 46.180 27.025 46.350 30.065 ;
        RECT 47.470 27.025 47.640 30.065 ;
        RECT 48.760 27.025 48.930 30.065 ;
        RECT 50.050 27.025 50.220 30.065 ;
        RECT 51.340 27.025 51.510 30.065 ;
        RECT 52.630 27.025 52.800 30.065 ;
        RECT 53.920 27.025 54.090 30.065 ;
        RECT 55.210 27.025 55.380 30.065 ;
        RECT 56.500 27.025 56.670 30.065 ;
        RECT 57.070 29.995 57.240 30.745 ;
        RECT 58.935 30.745 67.985 30.915 ;
        RECT 58.935 29.995 59.105 30.745 ;
        RECT 61.025 30.235 62.025 30.405 ;
        RECT 62.315 30.235 63.315 30.405 ;
        RECT 63.605 30.235 64.605 30.405 ;
        RECT 64.895 30.235 65.895 30.405 ;
        RECT 57.055 27.095 57.255 29.995 ;
        RECT 58.905 27.095 59.105 29.995 ;
        RECT 46.410 26.685 47.410 26.855 ;
        RECT 55.440 26.685 56.440 26.855 ;
        RECT 57.070 26.345 57.240 27.095 ;
        RECT 45.610 26.175 57.240 26.345 ;
        RECT 58.935 26.345 59.105 27.095 ;
        RECT 59.505 27.025 59.675 30.065 ;
        RECT 60.795 27.025 60.965 30.065 ;
        RECT 62.085 27.025 62.255 30.065 ;
        RECT 63.375 27.025 63.545 30.065 ;
        RECT 64.665 27.025 64.835 30.065 ;
        RECT 65.955 27.025 66.125 30.065 ;
        RECT 67.245 27.025 67.415 30.065 ;
        RECT 67.815 29.995 67.985 30.745 ;
        RECT 69.685 30.745 81.315 30.915 ;
        RECT 69.685 29.995 69.855 30.745 ;
        RECT 71.775 30.235 72.775 30.405 ;
        RECT 73.065 30.235 74.065 30.405 ;
        RECT 74.355 30.235 75.355 30.405 ;
        RECT 75.645 30.235 76.645 30.405 ;
        RECT 76.935 30.235 77.935 30.405 ;
        RECT 78.225 30.235 79.225 30.405 ;
        RECT 67.805 27.095 68.005 29.995 ;
        RECT 69.655 27.095 69.855 29.995 ;
        RECT 59.735 26.685 60.735 26.855 ;
        RECT 66.185 26.685 67.185 26.855 ;
        RECT 67.815 26.345 67.985 27.095 ;
        RECT 58.935 26.175 67.985 26.345 ;
        RECT 69.685 26.345 69.855 27.095 ;
        RECT 70.255 27.025 70.425 30.065 ;
        RECT 71.545 27.025 71.715 30.065 ;
        RECT 74.125 27.025 74.295 30.065 ;
        RECT 76.705 27.025 76.875 30.065 ;
        RECT 79.285 27.025 79.455 30.065 ;
        RECT 80.575 27.025 80.745 30.065 ;
        RECT 81.145 29.995 81.315 30.745 ;
        RECT 83.010 30.745 94.640 30.915 ;
        RECT 83.010 29.995 83.180 30.745 ;
        RECT 85.100 30.235 86.100 30.405 ;
        RECT 86.390 30.235 87.390 30.405 ;
        RECT 87.680 30.235 88.680 30.405 ;
        RECT 88.970 30.235 89.970 30.405 ;
        RECT 90.260 30.235 91.260 30.405 ;
        RECT 91.550 30.235 92.550 30.405 ;
        RECT 81.130 27.095 81.330 29.995 ;
        RECT 82.980 27.095 83.180 29.995 ;
        RECT 70.485 26.685 71.485 26.855 ;
        RECT 79.515 26.685 80.515 26.855 ;
        RECT 81.145 26.345 81.315 27.095 ;
        RECT 69.685 26.175 81.315 26.345 ;
        RECT 83.010 26.345 83.180 27.095 ;
        RECT 83.580 27.025 83.750 30.065 ;
        RECT 84.870 27.025 85.040 30.065 ;
        RECT 87.450 27.025 87.620 30.065 ;
        RECT 90.030 27.025 90.200 30.065 ;
        RECT 92.610 27.025 92.780 30.065 ;
        RECT 93.900 27.025 94.070 30.065 ;
        RECT 94.470 29.995 94.640 30.745 ;
        RECT 96.335 30.745 107.965 30.915 ;
        RECT 96.335 29.995 96.505 30.745 ;
        RECT 98.425 30.235 99.425 30.405 ;
        RECT 99.715 30.235 100.715 30.405 ;
        RECT 101.005 30.235 102.005 30.405 ;
        RECT 102.295 30.235 103.295 30.405 ;
        RECT 103.585 30.235 104.585 30.405 ;
        RECT 104.875 30.235 105.875 30.405 ;
        RECT 94.455 27.095 94.655 29.995 ;
        RECT 96.305 27.095 96.505 29.995 ;
        RECT 83.810 26.685 84.810 26.855 ;
        RECT 92.840 26.685 93.840 26.855 ;
        RECT 94.470 26.345 94.640 27.095 ;
        RECT 83.010 26.175 94.640 26.345 ;
        RECT 96.335 26.345 96.505 27.095 ;
        RECT 96.905 27.025 97.075 30.065 ;
        RECT 98.195 27.025 98.365 30.065 ;
        RECT 100.775 27.025 100.945 30.065 ;
        RECT 103.355 27.025 103.525 30.065 ;
        RECT 105.935 27.025 106.105 30.065 ;
        RECT 107.225 27.025 107.395 30.065 ;
        RECT 107.795 29.995 107.965 30.745 ;
        RECT 109.660 30.745 121.290 30.915 ;
        RECT 109.660 29.995 109.830 30.745 ;
        RECT 111.750 30.235 112.750 30.405 ;
        RECT 113.040 30.235 114.040 30.405 ;
        RECT 114.330 30.235 115.330 30.405 ;
        RECT 115.620 30.235 116.620 30.405 ;
        RECT 116.910 30.235 117.910 30.405 ;
        RECT 118.200 30.235 119.200 30.405 ;
        RECT 107.780 27.095 107.980 29.995 ;
        RECT 109.630 27.095 109.830 29.995 ;
        RECT 97.135 26.685 98.135 26.855 ;
        RECT 106.165 26.685 107.165 26.855 ;
        RECT 107.795 26.345 107.965 27.095 ;
        RECT 96.335 26.175 107.965 26.345 ;
        RECT 109.660 26.345 109.830 27.095 ;
        RECT 110.230 27.025 110.400 30.065 ;
        RECT 111.520 27.025 111.690 30.065 ;
        RECT 114.100 27.025 114.270 30.065 ;
        RECT 116.680 27.025 116.850 30.065 ;
        RECT 119.260 27.025 119.430 30.065 ;
        RECT 120.550 27.025 120.720 30.065 ;
        RECT 121.120 29.995 121.290 30.745 ;
        RECT 122.985 30.745 134.615 30.915 ;
        RECT 122.985 29.995 123.155 30.745 ;
        RECT 125.075 30.235 126.075 30.405 ;
        RECT 126.365 30.235 127.365 30.405 ;
        RECT 127.655 30.235 128.655 30.405 ;
        RECT 128.945 30.235 129.945 30.405 ;
        RECT 130.235 30.235 131.235 30.405 ;
        RECT 131.525 30.235 132.525 30.405 ;
        RECT 121.105 27.095 121.305 29.995 ;
        RECT 122.955 27.095 123.155 29.995 ;
        RECT 110.460 26.685 111.460 26.855 ;
        RECT 119.490 26.685 120.490 26.855 ;
        RECT 121.120 26.345 121.290 27.095 ;
        RECT 109.660 26.175 121.290 26.345 ;
        RECT 122.985 26.345 123.155 27.095 ;
        RECT 123.555 27.025 123.725 30.065 ;
        RECT 124.845 27.025 125.015 30.065 ;
        RECT 126.135 27.025 126.305 30.065 ;
        RECT 127.425 27.025 127.595 30.065 ;
        RECT 128.715 27.025 128.885 30.065 ;
        RECT 130.005 27.025 130.175 30.065 ;
        RECT 131.295 27.025 131.465 30.065 ;
        RECT 132.585 27.025 132.755 30.065 ;
        RECT 133.875 27.025 134.045 30.065 ;
        RECT 134.445 29.995 134.615 30.745 ;
        RECT 136.310 30.745 145.360 30.915 ;
        RECT 136.310 29.995 136.480 30.745 ;
        RECT 138.400 30.235 139.400 30.405 ;
        RECT 139.690 30.235 140.690 30.405 ;
        RECT 140.980 30.235 141.980 30.405 ;
        RECT 142.270 30.235 143.270 30.405 ;
        RECT 134.430 27.095 134.630 29.995 ;
        RECT 136.280 27.095 136.480 29.995 ;
        RECT 123.785 26.685 124.785 26.855 ;
        RECT 132.815 26.685 133.815 26.855 ;
        RECT 134.445 26.345 134.615 27.095 ;
        RECT 122.985 26.175 134.615 26.345 ;
        RECT 136.310 26.345 136.480 27.095 ;
        RECT 136.880 27.025 137.050 30.065 ;
        RECT 138.170 27.025 138.340 30.065 ;
        RECT 139.460 27.025 139.630 30.065 ;
        RECT 140.750 27.025 140.920 30.065 ;
        RECT 142.040 27.025 142.210 30.065 ;
        RECT 143.330 27.025 143.500 30.065 ;
        RECT 144.620 27.025 144.790 30.065 ;
        RECT 145.190 29.995 145.360 30.745 ;
        RECT 147.060 30.745 158.690 30.915 ;
        RECT 147.060 29.995 147.230 30.745 ;
        RECT 145.180 27.095 145.380 29.995 ;
        RECT 147.030 27.095 147.230 29.995 ;
        RECT 137.110 26.685 138.110 26.855 ;
        RECT 143.560 26.685 144.560 26.855 ;
        RECT 145.190 26.345 145.360 27.095 ;
        RECT 136.310 26.175 145.360 26.345 ;
        RECT 147.060 26.345 147.230 27.095 ;
        RECT 147.630 27.025 147.800 30.065 ;
        RECT 148.920 27.025 149.090 30.065 ;
        RECT 150.210 27.025 150.380 30.065 ;
        RECT 151.500 27.025 151.670 30.065 ;
        RECT 152.790 27.025 152.960 30.065 ;
        RECT 154.080 27.025 154.250 30.065 ;
        RECT 155.370 27.025 155.540 30.065 ;
        RECT 156.660 27.025 156.830 30.065 ;
        RECT 157.950 27.025 158.120 30.065 ;
        RECT 158.520 29.995 158.690 30.745 ;
        RECT 160.385 30.745 172.015 30.915 ;
        RECT 160.385 29.995 160.555 30.745 ;
        RECT 158.505 27.095 158.705 29.995 ;
        RECT 160.355 27.095 160.555 29.995 ;
        RECT 147.860 26.685 148.860 26.855 ;
        RECT 156.890 26.685 157.890 26.855 ;
        RECT 158.520 26.345 158.690 27.095 ;
        RECT 147.060 26.175 158.690 26.345 ;
        RECT 160.385 26.345 160.555 27.095 ;
        RECT 160.955 27.025 161.125 30.065 ;
        RECT 162.245 27.025 162.415 30.065 ;
        RECT 163.535 27.025 163.705 30.065 ;
        RECT 164.825 27.025 164.995 30.065 ;
        RECT 166.115 27.025 166.285 30.065 ;
        RECT 167.405 27.025 167.575 30.065 ;
        RECT 168.695 27.025 168.865 30.065 ;
        RECT 169.985 27.025 170.155 30.065 ;
        RECT 171.275 27.025 171.445 30.065 ;
        RECT 171.845 29.995 172.015 30.745 ;
        RECT 171.830 27.095 172.030 29.995 ;
        RECT 161.185 26.685 162.185 26.855 ;
        RECT 170.215 26.685 171.215 26.855 ;
        RECT 171.845 26.345 172.015 27.095 ;
        RECT 160.385 26.175 172.015 26.345 ;
        RECT 43.205 23.220 158.565 23.390 ;
        RECT 43.205 19.975 43.375 23.220 ;
        RECT 44.685 20.580 45.035 22.740 ;
        RECT 45.515 20.580 45.865 22.740 ;
        RECT 46.345 20.580 46.695 22.740 ;
        RECT 47.175 20.580 47.525 22.740 ;
        RECT 48.005 20.580 48.355 22.740 ;
        RECT 48.835 20.580 49.185 22.740 ;
        RECT 49.665 20.580 50.015 22.740 ;
        RECT 50.495 20.580 50.845 22.740 ;
        RECT 51.325 20.580 51.675 22.740 ;
        RECT 52.155 20.580 52.505 22.740 ;
        RECT 52.985 20.580 53.335 22.740 ;
        RECT 53.815 20.580 54.165 22.740 ;
        RECT 54.645 20.580 54.995 22.740 ;
        RECT 55.475 20.580 55.825 22.740 ;
        RECT 56.305 20.580 56.655 22.740 ;
        RECT 57.135 20.580 57.485 22.740 ;
        RECT 57.965 20.580 58.315 22.740 ;
        RECT 58.795 20.580 59.145 22.740 ;
        RECT 59.625 20.580 59.975 22.740 ;
        RECT 60.455 20.580 60.805 22.740 ;
        RECT 61.285 20.580 61.635 22.740 ;
        RECT 62.115 20.580 62.465 22.740 ;
        RECT 62.945 20.580 63.295 22.740 ;
        RECT 63.775 20.580 64.125 22.740 ;
        RECT 64.605 20.580 64.955 22.740 ;
        RECT 65.435 20.580 65.785 22.740 ;
        RECT 66.265 20.580 66.615 22.740 ;
        RECT 67.095 20.580 67.445 22.740 ;
        RECT 67.925 20.580 68.275 22.740 ;
        RECT 68.755 20.580 69.105 22.740 ;
        RECT 69.585 20.580 69.935 22.740 ;
        RECT 70.415 20.580 70.765 22.740 ;
        RECT 71.245 20.580 71.595 22.740 ;
        RECT 72.075 20.580 72.425 22.740 ;
        RECT 72.905 20.580 73.255 22.740 ;
        RECT 73.735 20.580 74.085 22.740 ;
        RECT 74.565 20.580 74.915 22.740 ;
        RECT 75.395 20.580 75.745 22.740 ;
        RECT 76.225 20.580 76.575 22.740 ;
        RECT 77.055 20.580 77.405 22.740 ;
        RECT 77.885 20.580 78.235 22.740 ;
        RECT 78.715 20.580 79.065 22.740 ;
        RECT 79.545 20.580 79.895 22.740 ;
        RECT 80.375 20.580 80.725 22.740 ;
        RECT 81.205 20.580 81.555 22.740 ;
        RECT 82.035 20.580 82.385 22.740 ;
        RECT 82.865 20.580 83.215 22.740 ;
        RECT 83.695 20.580 84.045 22.740 ;
        RECT 84.525 20.580 84.875 22.740 ;
        RECT 85.355 20.580 85.705 22.740 ;
        RECT 86.185 20.580 86.535 22.740 ;
        RECT 87.015 20.580 87.365 22.740 ;
        RECT 87.845 20.580 88.195 22.740 ;
        RECT 88.675 20.580 89.025 22.740 ;
        RECT 89.505 20.580 89.855 22.740 ;
        RECT 90.335 20.580 90.685 22.740 ;
        RECT 91.165 20.580 91.515 22.740 ;
        RECT 91.995 20.580 92.345 22.740 ;
        RECT 92.825 20.580 93.175 22.740 ;
        RECT 93.655 20.580 94.005 22.740 ;
        RECT 94.485 20.580 94.835 22.740 ;
        RECT 95.315 20.580 95.665 22.740 ;
        RECT 96.145 20.580 96.495 22.740 ;
        RECT 96.975 20.580 97.325 22.740 ;
        RECT 97.805 20.580 98.155 22.740 ;
        RECT 98.635 20.580 98.985 22.740 ;
        RECT 99.465 20.580 99.815 22.740 ;
        RECT 100.295 20.580 100.645 22.740 ;
        RECT 101.125 20.580 101.475 22.740 ;
        RECT 101.955 20.580 102.305 22.740 ;
        RECT 102.785 20.580 103.135 22.740 ;
        RECT 103.615 20.580 103.965 22.740 ;
        RECT 104.445 20.580 104.795 22.740 ;
        RECT 105.275 20.580 105.625 22.740 ;
        RECT 106.105 20.580 106.455 22.740 ;
        RECT 106.935 20.580 107.285 22.740 ;
        RECT 107.765 20.580 108.115 22.740 ;
        RECT 108.595 20.580 108.945 22.740 ;
        RECT 109.425 20.580 109.775 22.740 ;
        RECT 110.255 20.580 110.605 22.740 ;
        RECT 111.085 20.580 111.435 22.740 ;
        RECT 111.915 20.580 112.265 22.740 ;
        RECT 112.745 20.580 113.095 22.740 ;
        RECT 113.575 20.580 113.925 22.740 ;
        RECT 114.405 20.580 114.755 22.740 ;
        RECT 115.235 20.580 115.585 22.740 ;
        RECT 116.065 20.580 116.415 22.740 ;
        RECT 116.895 20.580 117.245 22.740 ;
        RECT 117.725 20.580 118.075 22.740 ;
        RECT 118.555 20.580 118.905 22.740 ;
        RECT 119.385 20.580 119.735 22.740 ;
        RECT 120.215 20.580 120.565 22.740 ;
        RECT 121.045 20.580 121.395 22.740 ;
        RECT 121.875 20.580 122.225 22.740 ;
        RECT 122.705 20.580 123.055 22.740 ;
        RECT 123.535 20.580 123.885 22.740 ;
        RECT 124.365 20.580 124.715 22.740 ;
        RECT 125.195 20.580 125.545 22.740 ;
        RECT 126.025 20.580 126.375 22.740 ;
        RECT 126.855 20.580 127.205 22.740 ;
        RECT 127.685 20.580 128.035 22.740 ;
        RECT 128.515 20.580 128.865 22.740 ;
        RECT 129.345 20.580 129.695 22.740 ;
        RECT 130.175 20.580 130.525 22.740 ;
        RECT 131.005 20.580 131.355 22.740 ;
        RECT 131.835 20.580 132.185 22.740 ;
        RECT 132.665 20.580 133.015 22.740 ;
        RECT 133.495 20.580 133.845 22.740 ;
        RECT 134.325 20.580 134.675 22.740 ;
        RECT 135.155 20.580 135.505 22.740 ;
        RECT 135.985 20.580 136.335 22.740 ;
        RECT 136.815 20.580 137.165 22.740 ;
        RECT 137.645 20.580 137.995 22.740 ;
        RECT 138.475 20.580 138.825 22.740 ;
        RECT 139.305 20.580 139.655 22.740 ;
        RECT 140.135 20.580 140.485 22.740 ;
        RECT 140.965 20.580 141.315 22.740 ;
        RECT 141.795 20.580 142.145 22.740 ;
        RECT 142.625 20.580 142.975 22.740 ;
        RECT 143.455 20.580 143.805 22.740 ;
        RECT 144.285 20.580 144.635 22.740 ;
        RECT 145.115 20.580 145.465 22.740 ;
        RECT 145.945 20.580 146.295 22.740 ;
        RECT 146.775 20.580 147.125 22.740 ;
        RECT 147.605 20.580 147.955 22.740 ;
        RECT 148.435 20.580 148.785 22.740 ;
        RECT 149.265 20.580 149.615 22.740 ;
        RECT 150.095 20.580 150.445 22.740 ;
        RECT 150.925 20.580 151.275 22.740 ;
        RECT 151.755 20.580 152.105 22.740 ;
        RECT 152.585 20.580 152.935 22.740 ;
        RECT 153.415 20.580 153.765 22.740 ;
        RECT 154.245 20.580 154.595 22.740 ;
        RECT 155.075 20.580 155.425 22.740 ;
        RECT 155.905 20.580 156.255 22.740 ;
        RECT 156.735 20.580 157.085 22.740 ;
        RECT 43.025 19.350 43.550 19.975 ;
        RECT 43.205 16.100 43.375 19.350 ;
        RECT 43.855 16.580 44.205 18.740 ;
        RECT 44.685 16.580 45.035 18.740 ;
        RECT 45.515 16.580 45.865 18.740 ;
        RECT 46.345 16.580 46.695 18.740 ;
        RECT 47.175 16.580 47.525 18.740 ;
        RECT 48.005 16.580 48.355 18.740 ;
        RECT 48.835 16.580 49.185 18.740 ;
        RECT 49.665 16.580 50.015 18.740 ;
        RECT 50.495 16.580 50.845 18.740 ;
        RECT 51.325 16.580 51.675 18.740 ;
        RECT 52.155 16.580 52.505 18.740 ;
        RECT 52.985 16.580 53.335 18.740 ;
        RECT 53.815 16.580 54.165 18.740 ;
        RECT 54.645 16.580 54.995 18.740 ;
        RECT 55.475 16.580 55.825 18.740 ;
        RECT 56.305 16.580 56.655 18.740 ;
        RECT 57.135 16.580 57.485 18.740 ;
        RECT 57.965 16.580 58.315 18.740 ;
        RECT 58.795 16.580 59.145 18.740 ;
        RECT 59.625 16.580 59.975 18.740 ;
        RECT 60.455 16.580 60.805 18.740 ;
        RECT 61.285 16.580 61.635 18.740 ;
        RECT 62.115 16.580 62.465 18.740 ;
        RECT 62.945 16.580 63.295 18.740 ;
        RECT 63.775 16.580 64.125 18.740 ;
        RECT 64.605 16.580 64.955 18.740 ;
        RECT 65.435 16.580 65.785 18.740 ;
        RECT 66.265 16.580 66.615 18.740 ;
        RECT 67.095 16.580 67.445 18.740 ;
        RECT 67.925 16.580 68.275 18.740 ;
        RECT 68.755 16.580 69.105 18.740 ;
        RECT 69.585 16.580 69.935 18.740 ;
        RECT 70.415 16.580 70.765 18.740 ;
        RECT 71.245 16.580 71.595 18.740 ;
        RECT 72.075 16.580 72.425 18.740 ;
        RECT 72.905 16.580 73.255 18.740 ;
        RECT 73.735 16.580 74.085 18.740 ;
        RECT 74.565 16.580 74.915 18.740 ;
        RECT 75.395 16.580 75.745 18.740 ;
        RECT 76.225 16.580 76.575 18.740 ;
        RECT 77.055 16.580 77.405 18.740 ;
        RECT 77.885 16.580 78.235 18.740 ;
        RECT 78.715 16.580 79.065 18.740 ;
        RECT 79.545 16.580 79.895 18.740 ;
        RECT 80.375 16.580 80.725 18.740 ;
        RECT 81.205 16.580 81.555 18.740 ;
        RECT 82.035 16.580 82.385 18.740 ;
        RECT 82.865 16.580 83.215 18.740 ;
        RECT 83.695 16.580 84.045 18.740 ;
        RECT 84.525 16.580 84.875 18.740 ;
        RECT 85.355 16.580 85.705 18.740 ;
        RECT 86.185 16.580 86.535 18.740 ;
        RECT 87.015 16.580 87.365 18.740 ;
        RECT 87.845 16.580 88.195 18.740 ;
        RECT 88.675 16.580 89.025 18.740 ;
        RECT 89.505 16.580 89.855 18.740 ;
        RECT 90.335 16.580 90.685 18.740 ;
        RECT 91.165 16.580 91.515 18.740 ;
        RECT 91.995 16.580 92.345 18.740 ;
        RECT 92.825 16.580 93.175 18.740 ;
        RECT 93.655 16.580 94.005 18.740 ;
        RECT 94.485 16.580 94.835 18.740 ;
        RECT 95.315 16.580 95.665 18.740 ;
        RECT 96.145 16.580 96.495 18.740 ;
        RECT 96.975 16.580 97.325 18.740 ;
        RECT 97.805 16.580 98.155 18.740 ;
        RECT 98.635 16.580 98.985 18.740 ;
        RECT 99.465 16.580 99.815 18.740 ;
        RECT 100.295 16.580 100.645 18.740 ;
        RECT 101.125 16.580 101.475 18.740 ;
        RECT 101.955 16.580 102.305 18.740 ;
        RECT 102.785 16.580 103.135 18.740 ;
        RECT 103.615 16.580 103.965 18.740 ;
        RECT 104.445 16.580 104.795 18.740 ;
        RECT 105.275 16.580 105.625 18.740 ;
        RECT 106.105 16.580 106.455 18.740 ;
        RECT 106.935 16.580 107.285 18.740 ;
        RECT 107.765 16.580 108.115 18.740 ;
        RECT 108.595 16.580 108.945 18.740 ;
        RECT 109.425 16.580 109.775 18.740 ;
        RECT 110.255 16.580 110.605 18.740 ;
        RECT 111.085 16.580 111.435 18.740 ;
        RECT 111.915 16.580 112.265 18.740 ;
        RECT 112.745 16.580 113.095 18.740 ;
        RECT 113.575 16.580 113.925 18.740 ;
        RECT 114.405 16.580 114.755 18.740 ;
        RECT 115.235 16.580 115.585 18.740 ;
        RECT 116.065 16.580 116.415 18.740 ;
        RECT 116.895 16.580 117.245 18.740 ;
        RECT 117.725 16.580 118.075 18.740 ;
        RECT 118.555 16.580 118.905 18.740 ;
        RECT 119.385 16.580 119.735 18.740 ;
        RECT 120.215 16.580 120.565 18.740 ;
        RECT 121.045 16.580 121.395 18.740 ;
        RECT 121.875 16.580 122.225 18.740 ;
        RECT 122.705 16.580 123.055 18.740 ;
        RECT 123.535 16.580 123.885 18.740 ;
        RECT 124.365 16.580 124.715 18.740 ;
        RECT 125.195 16.580 125.545 18.740 ;
        RECT 126.025 16.580 126.375 18.740 ;
        RECT 126.855 16.580 127.205 18.740 ;
        RECT 127.685 16.580 128.035 18.740 ;
        RECT 128.515 16.580 128.865 18.740 ;
        RECT 129.345 16.580 129.695 18.740 ;
        RECT 130.175 16.580 130.525 18.740 ;
        RECT 131.005 16.580 131.355 18.740 ;
        RECT 131.835 16.580 132.185 18.740 ;
        RECT 132.665 16.580 133.015 18.740 ;
        RECT 133.495 16.580 133.845 18.740 ;
        RECT 134.325 16.580 134.675 18.740 ;
        RECT 135.155 16.580 135.505 18.740 ;
        RECT 135.985 16.580 136.335 18.740 ;
        RECT 136.815 16.580 137.165 18.740 ;
        RECT 137.645 16.580 137.995 18.740 ;
        RECT 138.475 16.580 138.825 18.740 ;
        RECT 139.305 16.580 139.655 18.740 ;
        RECT 140.135 16.580 140.485 18.740 ;
        RECT 140.965 16.580 141.315 18.740 ;
        RECT 141.795 16.580 142.145 18.740 ;
        RECT 142.625 16.580 142.975 18.740 ;
        RECT 143.455 16.580 143.805 18.740 ;
        RECT 144.285 16.580 144.635 18.740 ;
        RECT 145.115 16.580 145.465 18.740 ;
        RECT 145.945 16.580 146.295 18.740 ;
        RECT 146.775 16.580 147.125 18.740 ;
        RECT 147.605 16.580 147.955 18.740 ;
        RECT 148.435 16.580 148.785 18.740 ;
        RECT 149.265 16.580 149.615 18.740 ;
        RECT 150.095 16.580 150.445 18.740 ;
        RECT 150.925 16.580 151.275 18.740 ;
        RECT 151.755 16.580 152.105 18.740 ;
        RECT 152.585 16.580 152.935 18.740 ;
        RECT 153.415 16.580 153.765 18.740 ;
        RECT 154.245 16.580 154.595 18.740 ;
        RECT 155.075 16.580 155.425 18.740 ;
        RECT 155.905 16.580 156.255 18.740 ;
        RECT 156.735 16.580 157.085 18.740 ;
        RECT 157.565 16.580 157.915 18.740 ;
        RECT 158.395 16.100 158.565 23.220 ;
        RECT 43.205 15.930 158.565 16.100 ;
      LAYER met1 ;
        RECT 73.775 52.800 127.325 53.200 ;
        RECT 43.905 51.900 44.155 51.935 ;
        RECT 44.735 51.900 44.985 51.935 ;
        RECT 45.565 51.900 45.815 51.935 ;
        RECT 46.395 51.900 46.645 51.935 ;
        RECT 47.225 51.900 47.475 51.935 ;
        RECT 48.055 51.900 48.305 51.935 ;
        RECT 48.885 51.900 49.135 51.935 ;
        RECT 49.715 51.900 49.965 51.935 ;
        RECT 50.545 51.900 50.795 51.935 ;
        RECT 51.375 51.900 51.625 51.935 ;
        RECT 52.205 51.900 52.455 51.935 ;
        RECT 53.035 51.900 53.285 51.935 ;
        RECT 53.865 51.900 54.115 51.935 ;
        RECT 54.695 51.900 54.945 51.935 ;
        RECT 55.525 51.900 55.775 51.935 ;
        RECT 56.355 51.900 56.605 51.935 ;
        RECT 57.185 51.900 57.435 51.935 ;
        RECT 58.015 51.900 58.265 51.935 ;
        RECT 58.845 51.900 59.095 51.935 ;
        RECT 59.675 51.900 59.925 51.935 ;
        RECT 60.505 51.900 60.755 51.935 ;
        RECT 61.335 51.900 61.585 51.935 ;
        RECT 62.165 51.900 62.415 51.935 ;
        RECT 62.995 51.900 63.245 51.935 ;
        RECT 63.825 51.900 64.075 51.935 ;
        RECT 64.655 51.900 64.905 51.935 ;
        RECT 65.485 51.900 65.735 51.935 ;
        RECT 66.315 51.900 66.565 51.935 ;
        RECT 67.145 51.900 67.395 51.935 ;
        RECT 67.975 51.900 68.225 51.935 ;
        RECT 68.805 51.900 69.055 51.935 ;
        RECT 69.635 51.900 69.885 51.935 ;
        RECT 70.465 51.900 70.715 51.935 ;
        RECT 71.295 51.900 71.545 51.935 ;
        RECT 72.125 51.900 72.375 51.935 ;
        RECT 72.955 51.900 73.205 51.935 ;
        RECT 43.900 49.875 45.000 51.900 ;
        RECT 45.550 49.875 46.650 51.900 ;
        RECT 47.225 49.875 48.325 51.900 ;
        RECT 48.875 49.875 49.975 51.900 ;
        RECT 50.545 49.875 51.650 51.900 ;
        RECT 52.200 49.875 53.300 51.900 ;
        RECT 53.865 49.875 54.975 51.900 ;
        RECT 55.525 49.875 56.625 51.900 ;
        RECT 57.175 49.875 58.275 51.900 ;
        RECT 58.845 49.875 59.950 51.900 ;
        RECT 60.500 49.875 61.600 51.900 ;
        RECT 62.165 49.875 63.275 51.900 ;
        RECT 63.825 49.875 64.925 51.900 ;
        RECT 65.475 49.875 66.575 51.900 ;
        RECT 67.145 49.875 68.250 51.900 ;
        RECT 68.800 49.875 69.900 51.900 ;
        RECT 70.465 49.875 71.575 51.900 ;
        RECT 72.125 49.875 73.225 51.900 ;
        RECT 73.775 49.875 74.900 52.800 ;
        RECT 75.445 51.900 75.695 51.935 ;
        RECT 76.275 51.900 76.525 51.935 ;
        RECT 77.105 51.900 77.355 51.935 ;
        RECT 77.935 51.900 78.185 51.935 ;
        RECT 78.765 51.900 79.015 51.935 ;
        RECT 79.595 51.900 79.845 51.935 ;
        RECT 80.425 51.900 80.675 51.935 ;
        RECT 81.255 51.900 81.505 51.935 ;
        RECT 82.085 51.900 82.335 51.935 ;
        RECT 82.915 51.900 83.165 51.935 ;
        RECT 83.745 51.900 83.995 51.935 ;
        RECT 84.575 51.900 84.825 51.935 ;
        RECT 85.405 51.900 85.655 51.935 ;
        RECT 86.235 51.900 86.485 51.935 ;
        RECT 87.065 51.900 87.315 51.935 ;
        RECT 87.895 51.900 88.145 51.935 ;
        RECT 88.725 51.900 88.975 51.935 ;
        RECT 89.555 51.900 89.805 51.935 ;
        RECT 90.385 51.900 90.635 51.935 ;
        RECT 91.215 51.900 91.465 51.935 ;
        RECT 92.045 51.900 92.295 51.935 ;
        RECT 92.875 51.900 93.125 51.935 ;
        RECT 93.705 51.900 93.955 51.935 ;
        RECT 94.535 51.900 94.785 51.935 ;
        RECT 95.365 51.900 95.615 51.935 ;
        RECT 96.195 51.900 96.445 51.935 ;
        RECT 97.025 51.900 97.275 51.935 ;
        RECT 97.855 51.900 98.105 51.935 ;
        RECT 98.685 51.900 98.935 51.935 ;
        RECT 99.515 51.900 99.765 51.935 ;
        RECT 100.345 51.900 100.595 51.935 ;
        RECT 101.175 51.900 101.425 51.935 ;
        RECT 102.005 51.900 102.255 51.935 ;
        RECT 102.835 51.900 103.085 51.935 ;
        RECT 103.665 51.900 103.915 51.935 ;
        RECT 104.495 51.900 104.745 51.935 ;
        RECT 105.325 51.900 105.575 51.935 ;
        RECT 106.155 51.900 106.405 51.935 ;
        RECT 106.985 51.900 107.235 51.935 ;
        RECT 107.815 51.900 108.065 51.935 ;
        RECT 108.645 51.900 108.895 51.935 ;
        RECT 109.475 51.900 109.725 51.935 ;
        RECT 110.305 51.900 110.555 51.935 ;
        RECT 111.135 51.900 111.385 51.935 ;
        RECT 111.965 51.900 112.215 51.935 ;
        RECT 112.795 51.900 113.045 51.935 ;
        RECT 113.625 51.900 113.875 51.935 ;
        RECT 114.455 51.900 114.705 51.935 ;
        RECT 115.285 51.900 115.535 51.935 ;
        RECT 116.115 51.900 116.365 51.935 ;
        RECT 116.945 51.900 117.195 51.935 ;
        RECT 117.775 51.900 118.025 51.935 ;
        RECT 118.605 51.900 118.855 51.935 ;
        RECT 119.435 51.900 119.685 51.935 ;
        RECT 120.265 51.900 120.515 51.935 ;
        RECT 121.095 51.900 121.345 51.935 ;
        RECT 121.925 51.900 122.175 51.935 ;
        RECT 122.755 51.900 123.005 51.935 ;
        RECT 123.585 51.900 123.835 51.935 ;
        RECT 124.415 51.900 124.665 51.935 ;
        RECT 125.245 51.900 125.495 51.935 ;
        RECT 126.075 51.900 126.325 51.935 ;
        RECT 126.905 51.900 127.155 51.935 ;
        RECT 127.735 51.900 127.985 51.935 ;
        RECT 128.565 51.900 128.815 51.935 ;
        RECT 129.395 51.900 129.645 51.935 ;
        RECT 130.225 51.900 130.475 51.935 ;
        RECT 131.055 51.900 131.305 51.935 ;
        RECT 131.885 51.900 132.135 51.935 ;
        RECT 132.715 51.900 132.965 51.935 ;
        RECT 133.545 51.900 133.795 51.935 ;
        RECT 134.375 51.900 134.625 51.935 ;
        RECT 135.205 51.900 135.455 51.935 ;
        RECT 136.035 51.900 136.285 51.935 ;
        RECT 136.865 51.900 137.115 51.935 ;
        RECT 137.695 51.900 137.945 51.935 ;
        RECT 138.525 51.900 138.775 51.935 ;
        RECT 139.355 51.900 139.605 51.935 ;
        RECT 140.185 51.900 140.435 51.935 ;
        RECT 141.015 51.900 141.265 51.935 ;
        RECT 141.845 51.900 142.095 51.935 ;
        RECT 142.675 51.900 142.925 51.935 ;
        RECT 143.505 51.900 143.755 51.935 ;
        RECT 144.335 51.900 144.585 51.935 ;
        RECT 145.165 51.900 145.415 51.935 ;
        RECT 145.995 51.900 146.245 51.935 ;
        RECT 146.825 51.900 147.075 51.935 ;
        RECT 147.655 51.900 147.905 51.935 ;
        RECT 148.485 51.900 148.735 51.935 ;
        RECT 149.315 51.900 149.565 51.935 ;
        RECT 150.145 51.900 150.395 51.935 ;
        RECT 150.975 51.900 151.225 51.935 ;
        RECT 151.805 51.900 152.055 51.935 ;
        RECT 152.635 51.900 152.885 51.935 ;
        RECT 153.465 51.900 153.715 51.935 ;
        RECT 154.295 51.900 154.545 51.935 ;
        RECT 155.125 51.900 155.375 51.935 ;
        RECT 155.955 51.900 156.205 51.935 ;
        RECT 156.785 51.900 157.035 51.935 ;
        RECT 157.615 51.900 157.865 51.935 ;
        RECT 75.445 49.875 76.550 51.900 ;
        RECT 77.100 49.875 78.200 51.900 ;
        RECT 78.765 49.875 79.875 51.900 ;
        RECT 80.425 49.875 81.525 51.900 ;
        RECT 82.075 49.875 83.175 51.900 ;
        RECT 83.745 49.875 84.850 51.900 ;
        RECT 85.400 49.875 86.500 51.900 ;
        RECT 87.065 49.875 88.175 51.900 ;
        RECT 88.725 49.875 89.825 51.900 ;
        RECT 90.375 49.875 91.475 51.900 ;
        RECT 92.025 49.875 93.125 51.900 ;
        RECT 93.700 49.875 94.800 51.900 ;
        RECT 95.365 49.875 96.475 51.900 ;
        RECT 97.025 49.875 98.125 51.900 ;
        RECT 98.675 49.875 99.775 51.900 ;
        RECT 100.345 49.875 101.450 51.900 ;
        RECT 102.000 49.875 103.100 51.900 ;
        RECT 103.650 49.875 104.750 51.900 ;
        RECT 105.325 49.875 106.425 51.900 ;
        RECT 106.975 49.875 108.075 51.900 ;
        RECT 108.645 49.875 109.750 51.900 ;
        RECT 110.300 49.875 111.400 51.900 ;
        RECT 111.965 49.875 113.075 51.900 ;
        RECT 113.625 49.875 114.725 51.900 ;
        RECT 115.275 49.875 116.375 51.900 ;
        RECT 116.945 49.875 118.050 51.900 ;
        RECT 118.600 49.875 119.700 51.900 ;
        RECT 120.265 49.875 121.375 51.900 ;
        RECT 121.925 49.875 123.025 51.900 ;
        RECT 123.575 49.875 124.675 51.900 ;
        RECT 125.245 49.875 126.350 51.900 ;
        RECT 126.900 49.875 128.000 51.900 ;
        RECT 128.565 49.875 129.675 51.900 ;
        RECT 130.225 49.875 131.325 51.900 ;
        RECT 131.875 49.875 132.975 51.900 ;
        RECT 133.545 49.875 134.650 51.900 ;
        RECT 135.200 49.875 136.300 51.900 ;
        RECT 136.865 49.875 137.975 51.900 ;
        RECT 138.525 49.875 139.625 51.900 ;
        RECT 140.175 49.875 141.275 51.900 ;
        RECT 141.845 49.875 142.950 51.900 ;
        RECT 143.500 49.875 144.600 51.900 ;
        RECT 145.165 49.875 146.275 51.900 ;
        RECT 146.825 49.875 147.925 51.900 ;
        RECT 148.475 49.875 149.575 51.900 ;
        RECT 150.145 49.875 151.250 51.900 ;
        RECT 151.800 49.875 152.900 51.900 ;
        RECT 153.465 49.875 154.575 51.900 ;
        RECT 155.125 49.875 156.225 51.900 ;
        RECT 156.775 49.875 157.875 51.900 ;
        RECT 43.905 49.830 44.155 49.875 ;
        RECT 44.735 49.830 44.985 49.875 ;
        RECT 45.565 49.830 45.815 49.875 ;
        RECT 46.395 49.830 46.645 49.875 ;
        RECT 47.225 49.830 47.475 49.875 ;
        RECT 48.055 49.830 48.305 49.875 ;
        RECT 48.885 49.830 49.135 49.875 ;
        RECT 49.715 49.830 49.965 49.875 ;
        RECT 50.545 49.830 50.795 49.875 ;
        RECT 51.375 49.830 51.625 49.875 ;
        RECT 52.205 49.830 52.455 49.875 ;
        RECT 53.035 49.830 53.285 49.875 ;
        RECT 53.865 49.830 54.115 49.875 ;
        RECT 54.695 49.830 54.945 49.875 ;
        RECT 55.525 49.830 55.775 49.875 ;
        RECT 56.355 49.830 56.605 49.875 ;
        RECT 57.185 49.830 57.435 49.875 ;
        RECT 58.015 49.830 58.265 49.875 ;
        RECT 58.845 49.830 59.095 49.875 ;
        RECT 59.675 49.830 59.925 49.875 ;
        RECT 60.505 49.830 60.755 49.875 ;
        RECT 61.335 49.830 61.585 49.875 ;
        RECT 62.165 49.830 62.415 49.875 ;
        RECT 62.995 49.830 63.245 49.875 ;
        RECT 63.825 49.830 64.075 49.875 ;
        RECT 64.655 49.830 64.905 49.875 ;
        RECT 65.485 49.830 65.735 49.875 ;
        RECT 66.315 49.830 66.565 49.875 ;
        RECT 67.145 49.830 67.395 49.875 ;
        RECT 67.975 49.830 68.225 49.875 ;
        RECT 68.805 49.830 69.055 49.875 ;
        RECT 69.635 49.830 69.885 49.875 ;
        RECT 70.465 49.830 70.715 49.875 ;
        RECT 71.295 49.830 71.545 49.875 ;
        RECT 72.125 49.830 72.375 49.875 ;
        RECT 72.955 49.830 73.205 49.875 ;
        RECT 73.785 49.830 74.035 49.875 ;
        RECT 74.615 49.830 74.865 49.875 ;
        RECT 75.445 49.830 75.695 49.875 ;
        RECT 76.275 49.830 76.525 49.875 ;
        RECT 77.105 49.830 77.355 49.875 ;
        RECT 77.935 49.830 78.185 49.875 ;
        RECT 78.765 49.830 79.015 49.875 ;
        RECT 79.595 49.830 79.845 49.875 ;
        RECT 80.425 49.830 80.675 49.875 ;
        RECT 81.255 49.830 81.505 49.875 ;
        RECT 82.085 49.830 82.335 49.875 ;
        RECT 82.915 49.830 83.165 49.875 ;
        RECT 83.745 49.830 83.995 49.875 ;
        RECT 84.575 49.830 84.825 49.875 ;
        RECT 85.405 49.830 85.655 49.875 ;
        RECT 86.235 49.830 86.485 49.875 ;
        RECT 87.065 49.830 87.315 49.875 ;
        RECT 87.895 49.830 88.145 49.875 ;
        RECT 88.725 49.830 88.975 49.875 ;
        RECT 89.555 49.830 89.805 49.875 ;
        RECT 90.385 49.830 90.635 49.875 ;
        RECT 91.215 49.830 91.465 49.875 ;
        RECT 92.045 49.830 92.295 49.875 ;
        RECT 92.875 49.830 93.125 49.875 ;
        RECT 93.705 49.830 93.955 49.875 ;
        RECT 94.535 49.830 94.785 49.875 ;
        RECT 95.365 49.830 95.615 49.875 ;
        RECT 96.195 49.830 96.445 49.875 ;
        RECT 97.025 49.830 97.275 49.875 ;
        RECT 97.855 49.830 98.105 49.875 ;
        RECT 98.685 49.830 98.935 49.875 ;
        RECT 99.515 49.830 99.765 49.875 ;
        RECT 100.345 49.830 100.595 49.875 ;
        RECT 101.175 49.830 101.425 49.875 ;
        RECT 102.005 49.830 102.255 49.875 ;
        RECT 102.835 49.830 103.085 49.875 ;
        RECT 103.665 49.830 103.915 49.875 ;
        RECT 104.495 49.830 104.745 49.875 ;
        RECT 105.325 49.830 105.575 49.875 ;
        RECT 106.155 49.830 106.405 49.875 ;
        RECT 106.985 49.830 107.235 49.875 ;
        RECT 107.815 49.830 108.065 49.875 ;
        RECT 108.645 49.830 108.895 49.875 ;
        RECT 109.475 49.830 109.725 49.875 ;
        RECT 110.305 49.830 110.555 49.875 ;
        RECT 111.135 49.830 111.385 49.875 ;
        RECT 111.965 49.830 112.215 49.875 ;
        RECT 112.795 49.830 113.045 49.875 ;
        RECT 113.625 49.830 113.875 49.875 ;
        RECT 114.455 49.830 114.705 49.875 ;
        RECT 115.285 49.830 115.535 49.875 ;
        RECT 116.115 49.830 116.365 49.875 ;
        RECT 116.945 49.830 117.195 49.875 ;
        RECT 117.775 49.830 118.025 49.875 ;
        RECT 118.605 49.830 118.855 49.875 ;
        RECT 119.435 49.830 119.685 49.875 ;
        RECT 120.265 49.830 120.515 49.875 ;
        RECT 121.095 49.830 121.345 49.875 ;
        RECT 121.925 49.830 122.175 49.875 ;
        RECT 122.755 49.830 123.005 49.875 ;
        RECT 123.585 49.830 123.835 49.875 ;
        RECT 124.415 49.830 124.665 49.875 ;
        RECT 125.245 49.830 125.495 49.875 ;
        RECT 126.075 49.830 126.325 49.875 ;
        RECT 126.905 49.830 127.155 49.875 ;
        RECT 127.735 49.830 127.985 49.875 ;
        RECT 128.565 49.830 128.815 49.875 ;
        RECT 129.395 49.830 129.645 49.875 ;
        RECT 130.225 49.830 130.475 49.875 ;
        RECT 131.055 49.830 131.305 49.875 ;
        RECT 131.885 49.830 132.135 49.875 ;
        RECT 132.715 49.830 132.965 49.875 ;
        RECT 133.545 49.830 133.795 49.875 ;
        RECT 134.375 49.830 134.625 49.875 ;
        RECT 135.205 49.830 135.455 49.875 ;
        RECT 136.035 49.830 136.285 49.875 ;
        RECT 136.865 49.830 137.115 49.875 ;
        RECT 137.695 49.830 137.945 49.875 ;
        RECT 138.525 49.830 138.775 49.875 ;
        RECT 139.355 49.830 139.605 49.875 ;
        RECT 140.185 49.830 140.435 49.875 ;
        RECT 141.015 49.830 141.265 49.875 ;
        RECT 141.845 49.830 142.095 49.875 ;
        RECT 142.675 49.830 142.925 49.875 ;
        RECT 143.505 49.830 143.755 49.875 ;
        RECT 144.335 49.830 144.585 49.875 ;
        RECT 145.165 49.830 145.415 49.875 ;
        RECT 145.995 49.830 146.245 49.875 ;
        RECT 146.825 49.830 147.075 49.875 ;
        RECT 147.655 49.830 147.905 49.875 ;
        RECT 148.485 49.830 148.735 49.875 ;
        RECT 149.315 49.830 149.565 49.875 ;
        RECT 150.145 49.830 150.395 49.875 ;
        RECT 150.975 49.830 151.225 49.875 ;
        RECT 151.805 49.830 152.055 49.875 ;
        RECT 152.635 49.830 152.885 49.875 ;
        RECT 153.465 49.830 153.715 49.875 ;
        RECT 154.295 49.830 154.545 49.875 ;
        RECT 155.125 49.830 155.375 49.875 ;
        RECT 155.955 49.830 156.205 49.875 ;
        RECT 156.785 49.830 157.035 49.875 ;
        RECT 157.615 49.830 157.865 49.875 ;
        RECT 18.200 48.550 43.550 49.175 ;
        RECT 18.225 30.000 19.900 48.550 ;
        RECT 44.735 47.900 44.985 47.940 ;
        RECT 45.565 47.900 45.815 47.940 ;
        RECT 46.395 47.900 46.645 47.940 ;
        RECT 47.225 47.900 47.475 47.940 ;
        RECT 48.055 47.900 48.305 47.940 ;
        RECT 48.885 47.900 49.135 47.940 ;
        RECT 49.715 47.900 49.965 47.940 ;
        RECT 50.545 47.900 50.795 47.940 ;
        RECT 51.375 47.900 51.625 47.940 ;
        RECT 52.205 47.900 52.455 47.940 ;
        RECT 53.035 47.900 53.285 47.940 ;
        RECT 53.865 47.900 54.115 47.940 ;
        RECT 54.695 47.900 54.945 47.940 ;
        RECT 55.525 47.900 55.775 47.940 ;
        RECT 56.355 47.900 56.605 47.940 ;
        RECT 57.185 47.900 57.435 47.940 ;
        RECT 58.015 47.900 58.265 47.940 ;
        RECT 58.845 47.900 59.095 47.940 ;
        RECT 59.675 47.900 59.925 47.940 ;
        RECT 60.505 47.900 60.755 47.940 ;
        RECT 61.335 47.900 61.585 47.940 ;
        RECT 62.165 47.900 62.415 47.940 ;
        RECT 62.995 47.900 63.245 47.940 ;
        RECT 63.825 47.900 64.075 47.940 ;
        RECT 64.655 47.900 64.905 47.940 ;
        RECT 65.485 47.900 65.735 47.940 ;
        RECT 66.315 47.900 66.565 47.940 ;
        RECT 67.145 47.900 67.395 47.940 ;
        RECT 67.975 47.900 68.225 47.940 ;
        RECT 68.805 47.900 69.055 47.940 ;
        RECT 69.635 47.900 69.885 47.940 ;
        RECT 70.465 47.900 70.715 47.940 ;
        RECT 71.295 47.900 71.545 47.940 ;
        RECT 72.125 47.900 72.375 47.940 ;
        RECT 72.955 47.900 73.205 47.940 ;
        RECT 73.785 47.900 74.035 47.940 ;
        RECT 74.615 47.900 74.865 47.940 ;
        RECT 75.445 47.900 75.695 47.940 ;
        RECT 76.275 47.900 76.525 47.940 ;
        RECT 77.105 47.900 77.355 47.940 ;
        RECT 77.935 47.900 78.185 47.940 ;
        RECT 78.765 47.900 79.015 47.940 ;
        RECT 79.595 47.900 79.845 47.940 ;
        RECT 80.425 47.900 80.675 47.940 ;
        RECT 81.255 47.900 81.505 47.940 ;
        RECT 82.085 47.900 82.335 47.940 ;
        RECT 82.915 47.900 83.165 47.940 ;
        RECT 83.745 47.900 83.995 47.940 ;
        RECT 84.575 47.900 84.825 47.940 ;
        RECT 85.405 47.900 85.655 47.940 ;
        RECT 86.235 47.900 86.485 47.940 ;
        RECT 87.065 47.900 87.315 47.940 ;
        RECT 87.895 47.900 88.145 47.940 ;
        RECT 88.725 47.900 88.975 47.940 ;
        RECT 89.555 47.900 89.805 47.940 ;
        RECT 90.385 47.900 90.635 47.940 ;
        RECT 91.215 47.900 91.465 47.940 ;
        RECT 92.045 47.900 92.295 47.940 ;
        RECT 92.875 47.900 93.125 47.940 ;
        RECT 93.705 47.900 93.955 47.940 ;
        RECT 94.535 47.900 94.785 47.940 ;
        RECT 95.365 47.900 95.615 47.940 ;
        RECT 96.195 47.900 96.445 47.940 ;
        RECT 97.025 47.900 97.275 47.940 ;
        RECT 97.855 47.900 98.105 47.940 ;
        RECT 98.685 47.900 98.935 47.940 ;
        RECT 99.515 47.900 99.765 47.940 ;
        RECT 100.345 47.900 100.595 47.940 ;
        RECT 101.175 47.900 101.425 47.940 ;
        RECT 102.005 47.900 102.255 47.940 ;
        RECT 102.835 47.900 103.085 47.940 ;
        RECT 103.665 47.900 103.915 47.940 ;
        RECT 104.495 47.900 104.745 47.940 ;
        RECT 105.325 47.900 105.575 47.940 ;
        RECT 106.155 47.900 106.405 47.940 ;
        RECT 106.985 47.900 107.235 47.940 ;
        RECT 107.815 47.900 108.065 47.940 ;
        RECT 108.645 47.900 108.895 47.940 ;
        RECT 109.475 47.900 109.725 47.940 ;
        RECT 110.305 47.900 110.555 47.940 ;
        RECT 111.135 47.900 111.385 47.940 ;
        RECT 111.965 47.900 112.215 47.940 ;
        RECT 112.795 47.900 113.045 47.940 ;
        RECT 113.625 47.900 113.875 47.940 ;
        RECT 114.455 47.900 114.705 47.940 ;
        RECT 115.285 47.900 115.535 47.940 ;
        RECT 116.115 47.900 116.365 47.940 ;
        RECT 116.945 47.900 117.195 47.940 ;
        RECT 117.775 47.900 118.025 47.940 ;
        RECT 118.605 47.900 118.855 47.940 ;
        RECT 119.435 47.900 119.685 47.940 ;
        RECT 120.265 47.900 120.515 47.940 ;
        RECT 121.095 47.900 121.345 47.940 ;
        RECT 121.925 47.900 122.175 47.940 ;
        RECT 122.755 47.900 123.005 47.940 ;
        RECT 123.585 47.900 123.835 47.940 ;
        RECT 124.415 47.900 124.665 47.940 ;
        RECT 125.245 47.900 125.495 47.940 ;
        RECT 126.075 47.900 126.325 47.940 ;
        RECT 126.905 47.900 127.155 47.940 ;
        RECT 127.735 47.900 127.985 47.940 ;
        RECT 128.565 47.900 128.815 47.940 ;
        RECT 129.395 47.900 129.645 47.940 ;
        RECT 130.225 47.900 130.475 47.940 ;
        RECT 131.055 47.900 131.305 47.940 ;
        RECT 131.885 47.900 132.135 47.940 ;
        RECT 132.715 47.900 132.965 47.940 ;
        RECT 133.545 47.900 133.795 47.940 ;
        RECT 134.375 47.900 134.625 47.940 ;
        RECT 135.205 47.900 135.455 47.940 ;
        RECT 136.035 47.900 136.285 47.940 ;
        RECT 136.865 47.900 137.115 47.940 ;
        RECT 137.695 47.900 137.945 47.940 ;
        RECT 138.525 47.900 138.775 47.940 ;
        RECT 139.355 47.900 139.605 47.940 ;
        RECT 140.185 47.900 140.435 47.940 ;
        RECT 141.015 47.900 141.265 47.940 ;
        RECT 141.845 47.900 142.095 47.940 ;
        RECT 142.675 47.900 142.925 47.940 ;
        RECT 143.505 47.900 143.755 47.940 ;
        RECT 144.335 47.900 144.585 47.940 ;
        RECT 145.165 47.900 145.415 47.940 ;
        RECT 145.995 47.900 146.245 47.940 ;
        RECT 146.825 47.900 147.075 47.940 ;
        RECT 147.655 47.900 147.905 47.940 ;
        RECT 148.485 47.900 148.735 47.940 ;
        RECT 149.315 47.900 149.565 47.940 ;
        RECT 150.145 47.900 150.395 47.940 ;
        RECT 150.975 47.900 151.225 47.940 ;
        RECT 151.805 47.900 152.055 47.940 ;
        RECT 152.635 47.900 152.885 47.940 ;
        RECT 153.465 47.900 153.715 47.940 ;
        RECT 154.295 47.900 154.545 47.940 ;
        RECT 155.125 47.900 155.375 47.940 ;
        RECT 155.955 47.900 156.205 47.940 ;
        RECT 156.785 47.900 157.035 47.940 ;
        RECT 44.725 45.875 45.825 47.900 ;
        RECT 46.375 45.875 47.500 47.900 ;
        RECT 48.050 45.875 49.150 47.900 ;
        RECT 49.700 45.875 50.800 47.900 ;
        RECT 51.375 45.875 52.475 47.900 ;
        RECT 53.025 45.875 54.125 47.900 ;
        RECT 54.675 45.875 55.775 47.900 ;
        RECT 56.350 45.875 57.450 47.900 ;
        RECT 44.735 45.835 44.985 45.875 ;
        RECT 45.565 45.835 45.815 45.875 ;
        RECT 46.395 45.835 46.645 45.875 ;
        RECT 47.225 45.835 47.475 45.875 ;
        RECT 48.055 45.835 48.305 45.875 ;
        RECT 48.885 45.835 49.135 45.875 ;
        RECT 49.715 45.835 49.965 45.875 ;
        RECT 50.545 45.835 50.795 45.875 ;
        RECT 51.375 45.835 51.625 45.875 ;
        RECT 52.205 45.835 52.455 45.875 ;
        RECT 53.035 45.835 53.285 45.875 ;
        RECT 53.865 45.835 54.115 45.875 ;
        RECT 54.695 45.835 54.945 45.875 ;
        RECT 55.525 45.835 55.775 45.875 ;
        RECT 56.355 45.835 56.605 45.875 ;
        RECT 57.185 45.835 57.435 45.875 ;
        RECT 58.000 44.800 59.125 47.900 ;
        RECT 59.675 45.875 60.775 47.900 ;
        RECT 61.325 45.875 62.425 47.900 ;
        RECT 62.995 45.875 64.100 47.900 ;
        RECT 64.650 45.875 65.750 47.900 ;
        RECT 66.300 45.875 67.400 47.900 ;
        RECT 67.975 45.875 69.075 47.900 ;
        RECT 69.625 45.875 70.725 47.900 ;
        RECT 71.295 45.875 72.400 47.900 ;
        RECT 72.950 45.875 74.050 47.900 ;
        RECT 74.600 45.875 75.700 47.900 ;
        RECT 76.275 45.875 77.375 47.900 ;
        RECT 77.925 45.875 79.025 47.900 ;
        RECT 79.595 45.875 80.700 47.900 ;
        RECT 81.250 45.875 82.350 47.900 ;
        RECT 82.900 45.875 84.000 47.900 ;
        RECT 84.575 45.875 85.675 47.900 ;
        RECT 86.225 45.875 87.325 47.900 ;
        RECT 87.895 45.875 89.000 47.900 ;
        RECT 89.550 45.875 90.650 47.900 ;
        RECT 91.215 45.875 92.325 47.900 ;
        RECT 92.875 45.875 93.975 47.900 ;
        RECT 94.525 45.875 95.625 47.900 ;
        RECT 96.195 45.875 97.300 47.900 ;
        RECT 97.850 45.875 98.950 47.900 ;
        RECT 99.515 45.875 100.625 47.900 ;
        RECT 101.175 45.875 102.275 47.900 ;
        RECT 102.825 45.875 103.925 47.900 ;
        RECT 104.495 45.875 105.600 47.900 ;
        RECT 106.150 45.875 107.250 47.900 ;
        RECT 107.800 45.875 108.900 47.900 ;
        RECT 109.475 45.875 110.575 47.900 ;
        RECT 111.125 45.875 112.225 47.900 ;
        RECT 112.795 45.875 113.900 47.900 ;
        RECT 114.450 45.875 115.550 47.900 ;
        RECT 116.100 45.875 117.200 47.900 ;
        RECT 117.750 45.875 118.855 47.900 ;
        RECT 119.425 45.875 120.525 47.900 ;
        RECT 121.095 45.875 122.200 47.900 ;
        RECT 122.750 45.875 123.850 47.900 ;
        RECT 124.400 45.875 125.500 47.900 ;
        RECT 59.675 45.835 59.925 45.875 ;
        RECT 60.505 45.835 60.755 45.875 ;
        RECT 61.335 45.835 61.585 45.875 ;
        RECT 62.165 45.835 62.415 45.875 ;
        RECT 62.995 45.835 63.245 45.875 ;
        RECT 63.825 45.835 64.075 45.875 ;
        RECT 64.655 45.835 64.905 45.875 ;
        RECT 65.485 45.835 65.735 45.875 ;
        RECT 66.315 45.835 66.565 45.875 ;
        RECT 67.145 45.835 67.395 45.875 ;
        RECT 67.975 45.835 68.225 45.875 ;
        RECT 68.805 45.835 69.055 45.875 ;
        RECT 69.635 45.835 69.885 45.875 ;
        RECT 70.465 45.835 70.715 45.875 ;
        RECT 71.295 45.835 71.545 45.875 ;
        RECT 72.125 45.835 72.375 45.875 ;
        RECT 72.955 45.835 73.205 45.875 ;
        RECT 73.785 45.835 74.035 45.875 ;
        RECT 74.615 45.835 74.865 45.875 ;
        RECT 75.445 45.835 75.695 45.875 ;
        RECT 76.275 45.835 76.525 45.875 ;
        RECT 77.105 45.835 77.355 45.875 ;
        RECT 77.935 45.835 78.185 45.875 ;
        RECT 78.765 45.835 79.015 45.875 ;
        RECT 79.595 45.835 79.845 45.875 ;
        RECT 80.425 45.835 80.675 45.875 ;
        RECT 81.255 45.835 81.505 45.875 ;
        RECT 82.085 45.835 82.335 45.875 ;
        RECT 82.915 45.835 83.165 45.875 ;
        RECT 83.745 45.835 83.995 45.875 ;
        RECT 84.575 45.835 84.825 45.875 ;
        RECT 85.405 45.835 85.655 45.875 ;
        RECT 86.235 45.835 86.485 45.875 ;
        RECT 87.065 45.835 87.315 45.875 ;
        RECT 87.895 45.835 88.145 45.875 ;
        RECT 88.725 45.835 88.975 45.875 ;
        RECT 89.555 45.835 89.805 45.875 ;
        RECT 90.385 45.835 90.635 45.875 ;
        RECT 91.215 45.835 91.465 45.875 ;
        RECT 92.045 45.835 92.295 45.875 ;
        RECT 92.875 45.835 93.125 45.875 ;
        RECT 93.705 45.835 93.955 45.875 ;
        RECT 94.535 45.835 94.785 45.875 ;
        RECT 95.365 45.835 95.615 45.875 ;
        RECT 96.195 45.835 96.445 45.875 ;
        RECT 97.025 45.835 97.275 45.875 ;
        RECT 97.855 45.835 98.105 45.875 ;
        RECT 98.685 45.835 98.935 45.875 ;
        RECT 99.515 45.835 99.765 45.875 ;
        RECT 100.345 45.835 100.595 45.875 ;
        RECT 101.175 45.835 101.425 45.875 ;
        RECT 102.005 45.835 102.255 45.875 ;
        RECT 102.835 45.835 103.085 45.875 ;
        RECT 103.665 45.835 103.915 45.875 ;
        RECT 104.495 45.835 104.745 45.875 ;
        RECT 105.325 45.835 105.575 45.875 ;
        RECT 106.155 45.835 106.405 45.875 ;
        RECT 106.985 45.835 107.235 45.875 ;
        RECT 107.815 45.835 108.065 45.875 ;
        RECT 108.645 45.835 108.895 45.875 ;
        RECT 109.475 45.835 109.725 45.875 ;
        RECT 110.305 45.835 110.555 45.875 ;
        RECT 111.135 45.835 111.385 45.875 ;
        RECT 111.965 45.835 112.215 45.875 ;
        RECT 112.795 45.835 113.045 45.875 ;
        RECT 113.625 45.835 113.875 45.875 ;
        RECT 114.455 45.835 114.705 45.875 ;
        RECT 115.285 45.835 115.535 45.875 ;
        RECT 116.115 45.835 116.365 45.875 ;
        RECT 116.945 45.835 117.195 45.875 ;
        RECT 117.775 45.835 118.025 45.875 ;
        RECT 118.605 45.835 118.855 45.875 ;
        RECT 119.435 45.835 119.685 45.875 ;
        RECT 120.265 45.835 120.515 45.875 ;
        RECT 121.095 45.835 121.345 45.875 ;
        RECT 121.925 45.835 122.175 45.875 ;
        RECT 122.755 45.835 123.005 45.875 ;
        RECT 123.585 45.835 123.835 45.875 ;
        RECT 124.415 45.835 124.665 45.875 ;
        RECT 125.245 45.835 125.495 45.875 ;
        RECT 125.900 44.800 126.500 47.900 ;
        RECT 126.725 45.325 127.325 47.900 ;
        RECT 127.725 45.875 128.825 47.900 ;
        RECT 129.395 45.875 130.500 47.900 ;
        RECT 131.050 45.875 132.150 47.900 ;
        RECT 132.715 45.875 133.825 47.900 ;
        RECT 134.375 45.875 135.475 47.900 ;
        RECT 136.025 45.875 137.125 47.900 ;
        RECT 137.675 45.875 138.775 47.900 ;
        RECT 139.350 45.875 140.450 47.900 ;
        RECT 141.000 45.875 142.100 47.900 ;
        RECT 142.650 45.875 143.755 47.900 ;
        RECT 144.325 45.875 145.425 47.900 ;
        RECT 145.995 45.875 147.100 47.900 ;
        RECT 147.650 45.875 148.750 47.900 ;
        RECT 149.300 45.875 150.400 47.900 ;
        RECT 150.975 45.875 152.075 47.900 ;
        RECT 152.625 45.875 153.725 47.900 ;
        RECT 154.275 45.875 155.375 47.900 ;
        RECT 155.950 45.875 157.050 47.900 ;
        RECT 127.735 45.835 127.985 45.875 ;
        RECT 128.565 45.835 128.815 45.875 ;
        RECT 129.395 45.835 129.645 45.875 ;
        RECT 130.225 45.835 130.475 45.875 ;
        RECT 131.055 45.835 131.305 45.875 ;
        RECT 131.885 45.835 132.135 45.875 ;
        RECT 132.715 45.835 132.965 45.875 ;
        RECT 133.545 45.835 133.795 45.875 ;
        RECT 134.375 45.835 134.625 45.875 ;
        RECT 135.205 45.835 135.455 45.875 ;
        RECT 136.035 45.835 136.285 45.875 ;
        RECT 136.865 45.835 137.115 45.875 ;
        RECT 137.695 45.835 137.945 45.875 ;
        RECT 138.525 45.835 138.775 45.875 ;
        RECT 139.355 45.835 139.605 45.875 ;
        RECT 140.185 45.835 140.435 45.875 ;
        RECT 141.015 45.835 141.265 45.875 ;
        RECT 141.845 45.835 142.095 45.875 ;
        RECT 142.675 45.835 142.925 45.875 ;
        RECT 143.505 45.835 143.755 45.875 ;
        RECT 144.335 45.835 144.585 45.875 ;
        RECT 145.165 45.835 145.415 45.875 ;
        RECT 145.995 45.835 146.245 45.875 ;
        RECT 146.825 45.835 147.075 45.875 ;
        RECT 147.655 45.835 147.905 45.875 ;
        RECT 148.485 45.835 148.735 45.875 ;
        RECT 149.315 45.835 149.565 45.875 ;
        RECT 150.145 45.835 150.395 45.875 ;
        RECT 150.975 45.835 151.225 45.875 ;
        RECT 151.805 45.835 152.055 45.875 ;
        RECT 152.635 45.835 152.885 45.875 ;
        RECT 153.465 45.835 153.715 45.875 ;
        RECT 154.295 45.835 154.545 45.875 ;
        RECT 155.125 45.835 155.375 45.875 ;
        RECT 155.955 45.835 156.205 45.875 ;
        RECT 156.785 45.835 157.035 45.875 ;
        RECT 20.850 44.470 21.975 44.475 ;
        RECT 20.850 43.725 172.205 44.470 ;
        RECT 21.105 43.720 172.205 43.725 ;
        RECT 21.355 41.420 21.880 43.720 ;
        RECT 22.355 41.825 23.205 43.245 ;
        RECT 22.355 41.595 23.315 41.825 ;
        RECT 23.455 41.670 28.655 41.845 ;
        RECT 28.855 41.825 29.705 43.245 ;
        RECT 21.355 32.370 23.205 41.420 ;
        RECT 23.455 41.390 23.630 41.670 ;
        RECT 23.365 32.390 23.630 41.390 ;
        RECT 23.455 32.370 23.630 32.390 ;
        RECT 24.505 32.370 25.030 41.395 ;
        RECT 25.980 41.390 26.155 41.670 ;
        RECT 25.945 32.390 26.175 41.390 ;
        RECT 27.080 32.370 27.605 41.395 ;
        RECT 28.480 41.390 28.655 41.670 ;
        RECT 28.805 41.595 29.765 41.825 ;
        RECT 30.255 41.420 30.780 43.720 ;
        RECT 29.855 41.390 30.780 41.420 ;
        RECT 28.480 32.395 28.755 41.390 ;
        RECT 28.525 32.390 28.755 32.395 ;
        RECT 29.815 32.390 30.780 41.390 ;
        RECT 29.855 32.370 30.780 32.390 ;
        RECT 32.105 41.420 32.630 43.720 ;
        RECT 33.105 41.825 33.955 43.245 ;
        RECT 33.105 41.595 34.065 41.825 ;
        RECT 34.205 41.670 41.980 41.845 ;
        RECT 42.230 41.825 43.080 43.245 ;
        RECT 32.105 32.370 33.955 41.420 ;
        RECT 34.205 41.390 34.380 41.670 ;
        RECT 34.115 32.390 34.380 41.390 ;
        RECT 34.205 32.370 34.380 32.390 ;
        RECT 35.255 32.370 35.780 41.395 ;
        RECT 36.730 41.390 36.905 41.670 ;
        RECT 36.695 32.390 36.925 41.390 ;
        RECT 37.830 32.370 38.355 41.395 ;
        RECT 39.305 41.390 39.480 41.670 ;
        RECT 39.275 32.390 39.505 41.390 ;
        RECT 40.405 32.370 40.930 41.395 ;
        RECT 41.805 41.390 41.980 41.670 ;
        RECT 42.135 41.595 43.095 41.825 ;
        RECT 43.580 41.420 44.105 43.720 ;
        RECT 43.180 41.390 44.105 41.420 ;
        RECT 41.805 32.395 42.085 41.390 ;
        RECT 41.855 32.390 42.085 32.395 ;
        RECT 43.145 32.390 44.105 41.390 ;
        RECT 43.180 32.370 44.105 32.390 ;
        RECT 45.430 41.420 45.955 43.720 ;
        RECT 46.430 41.825 47.280 43.245 ;
        RECT 46.430 41.595 47.390 41.825 ;
        RECT 47.530 41.670 55.305 41.845 ;
        RECT 55.555 41.825 56.405 43.245 ;
        RECT 45.430 32.370 47.280 41.420 ;
        RECT 47.530 41.390 47.705 41.670 ;
        RECT 47.440 32.390 47.705 41.390 ;
        RECT 47.530 32.370 47.705 32.390 ;
        RECT 48.580 32.370 49.105 41.395 ;
        RECT 50.055 41.390 50.230 41.670 ;
        RECT 50.020 32.390 50.250 41.390 ;
        RECT 51.155 32.370 51.680 41.395 ;
        RECT 52.630 41.390 52.805 41.670 ;
        RECT 52.600 32.390 52.830 41.390 ;
        RECT 53.730 32.370 54.255 41.395 ;
        RECT 55.130 41.390 55.305 41.670 ;
        RECT 55.460 41.595 56.420 41.825 ;
        RECT 56.905 41.420 57.430 43.720 ;
        RECT 56.505 41.390 57.430 41.420 ;
        RECT 55.130 32.395 55.410 41.390 ;
        RECT 55.180 32.390 55.410 32.395 ;
        RECT 56.470 32.390 57.430 41.390 ;
        RECT 56.505 32.370 57.430 32.390 ;
        RECT 58.755 41.420 59.280 43.720 ;
        RECT 59.755 41.825 60.605 43.245 ;
        RECT 59.755 41.595 60.715 41.825 ;
        RECT 60.855 41.670 66.055 41.845 ;
        RECT 66.255 41.825 67.105 43.245 ;
        RECT 58.755 32.370 60.605 41.420 ;
        RECT 60.855 41.390 61.030 41.670 ;
        RECT 60.765 32.390 61.030 41.390 ;
        RECT 60.855 32.370 61.030 32.390 ;
        RECT 61.905 32.370 62.430 41.395 ;
        RECT 63.380 41.390 63.555 41.670 ;
        RECT 63.345 32.390 63.575 41.390 ;
        RECT 64.480 32.370 65.005 41.395 ;
        RECT 65.880 41.390 66.055 41.670 ;
        RECT 66.205 41.595 67.165 41.825 ;
        RECT 67.655 41.420 68.180 43.720 ;
        RECT 67.255 41.390 68.180 41.420 ;
        RECT 65.880 32.395 66.155 41.390 ;
        RECT 65.925 32.390 66.155 32.395 ;
        RECT 67.215 32.390 68.180 41.390 ;
        RECT 67.255 32.370 68.180 32.390 ;
        RECT 69.505 41.420 70.030 43.720 ;
        RECT 70.505 41.825 71.355 43.245 ;
        RECT 70.505 41.595 71.465 41.825 ;
        RECT 71.605 41.670 79.380 41.845 ;
        RECT 79.630 41.825 80.480 43.245 ;
        RECT 69.505 32.370 71.355 41.420 ;
        RECT 71.605 41.390 71.780 41.670 ;
        RECT 74.130 41.390 74.305 41.670 ;
        RECT 76.705 41.390 76.880 41.670 ;
        RECT 79.205 41.390 79.380 41.670 ;
        RECT 79.535 41.595 80.495 41.825 ;
        RECT 80.980 41.420 81.505 43.720 ;
        RECT 80.580 41.390 81.505 41.420 ;
        RECT 71.515 32.390 71.780 41.390 ;
        RECT 74.095 32.390 74.325 41.390 ;
        RECT 76.675 32.390 76.905 41.390 ;
        RECT 79.205 32.395 79.485 41.390 ;
        RECT 79.255 32.390 79.485 32.395 ;
        RECT 80.545 32.390 81.505 41.390 ;
        RECT 71.605 32.370 71.780 32.390 ;
        RECT 80.580 32.370 81.505 32.390 ;
        RECT 82.830 41.420 83.355 43.720 ;
        RECT 83.830 41.825 84.680 43.245 ;
        RECT 83.830 41.595 84.790 41.825 ;
        RECT 84.930 41.670 92.705 41.845 ;
        RECT 92.955 41.825 93.805 43.245 ;
        RECT 82.830 32.370 84.680 41.420 ;
        RECT 84.930 41.390 85.105 41.670 ;
        RECT 87.455 41.390 87.630 41.670 ;
        RECT 90.030 41.390 90.205 41.670 ;
        RECT 92.530 41.390 92.705 41.670 ;
        RECT 92.860 41.595 93.820 41.825 ;
        RECT 94.305 41.420 94.830 43.720 ;
        RECT 93.905 41.390 94.830 41.420 ;
        RECT 84.840 32.390 85.105 41.390 ;
        RECT 87.420 32.390 87.650 41.390 ;
        RECT 90.000 32.390 90.230 41.390 ;
        RECT 92.530 32.395 92.810 41.390 ;
        RECT 92.580 32.390 92.810 32.395 ;
        RECT 93.870 32.390 94.830 41.390 ;
        RECT 84.930 32.370 85.105 32.390 ;
        RECT 93.905 32.370 94.830 32.390 ;
        RECT 96.155 41.420 96.680 43.720 ;
        RECT 97.155 41.825 98.005 43.245 ;
        RECT 97.155 41.595 98.115 41.825 ;
        RECT 98.255 41.670 106.030 41.845 ;
        RECT 106.280 41.825 107.130 43.245 ;
        RECT 96.155 32.370 98.005 41.420 ;
        RECT 98.255 41.390 98.430 41.670 ;
        RECT 100.780 41.390 100.955 41.670 ;
        RECT 103.355 41.390 103.530 41.670 ;
        RECT 105.855 41.390 106.030 41.670 ;
        RECT 106.185 41.595 107.145 41.825 ;
        RECT 107.630 41.420 108.155 43.720 ;
        RECT 107.230 41.390 108.155 41.420 ;
        RECT 98.165 32.390 98.430 41.390 ;
        RECT 100.745 32.390 100.975 41.390 ;
        RECT 103.325 32.390 103.555 41.390 ;
        RECT 105.855 32.395 106.135 41.390 ;
        RECT 105.905 32.390 106.135 32.395 ;
        RECT 107.195 32.390 108.155 41.390 ;
        RECT 98.255 32.370 98.430 32.390 ;
        RECT 107.230 32.370 108.155 32.390 ;
        RECT 109.480 41.420 110.005 43.720 ;
        RECT 110.480 41.825 111.330 43.245 ;
        RECT 110.480 41.595 111.440 41.825 ;
        RECT 111.580 41.670 119.355 41.845 ;
        RECT 119.605 41.825 120.455 43.245 ;
        RECT 109.480 32.370 111.330 41.420 ;
        RECT 111.580 41.390 111.755 41.670 ;
        RECT 114.105 41.390 114.280 41.670 ;
        RECT 116.680 41.390 116.855 41.670 ;
        RECT 119.180 41.390 119.355 41.670 ;
        RECT 119.510 41.595 120.470 41.825 ;
        RECT 120.955 41.420 121.480 43.720 ;
        RECT 120.555 41.390 121.480 41.420 ;
        RECT 111.490 32.390 111.755 41.390 ;
        RECT 114.070 32.390 114.300 41.390 ;
        RECT 116.650 32.390 116.880 41.390 ;
        RECT 119.180 32.395 119.460 41.390 ;
        RECT 119.230 32.390 119.460 32.395 ;
        RECT 120.520 32.390 121.480 41.390 ;
        RECT 111.580 32.370 111.755 32.390 ;
        RECT 120.555 32.370 121.480 32.390 ;
        RECT 122.805 41.420 123.330 43.720 ;
        RECT 123.805 41.825 124.655 43.245 ;
        RECT 123.805 41.595 124.765 41.825 ;
        RECT 124.905 41.670 132.680 41.845 ;
        RECT 132.930 41.825 133.780 43.245 ;
        RECT 122.805 32.370 124.655 41.420 ;
        RECT 124.905 41.390 125.080 41.670 ;
        RECT 124.815 32.390 125.080 41.390 ;
        RECT 124.905 32.370 125.080 32.390 ;
        RECT 125.955 32.370 126.480 41.395 ;
        RECT 127.430 41.390 127.605 41.670 ;
        RECT 127.395 32.390 127.625 41.390 ;
        RECT 128.530 32.370 129.055 41.395 ;
        RECT 130.005 41.390 130.180 41.670 ;
        RECT 129.975 32.390 130.205 41.390 ;
        RECT 131.105 32.370 131.630 41.395 ;
        RECT 132.505 41.390 132.680 41.670 ;
        RECT 132.835 41.595 133.795 41.825 ;
        RECT 134.280 41.420 134.805 43.720 ;
        RECT 133.880 41.390 134.805 41.420 ;
        RECT 132.505 32.395 132.785 41.390 ;
        RECT 132.555 32.390 132.785 32.395 ;
        RECT 133.845 32.390 134.805 41.390 ;
        RECT 133.880 32.370 134.805 32.390 ;
        RECT 136.130 41.420 136.655 43.720 ;
        RECT 137.130 41.825 137.980 43.245 ;
        RECT 137.130 41.595 138.090 41.825 ;
        RECT 138.230 41.670 143.430 41.845 ;
        RECT 143.630 41.825 144.480 43.245 ;
        RECT 136.130 32.370 137.980 41.420 ;
        RECT 138.230 41.390 138.405 41.670 ;
        RECT 138.140 32.390 138.405 41.390 ;
        RECT 138.230 32.370 138.405 32.390 ;
        RECT 139.280 32.370 139.805 41.395 ;
        RECT 140.755 41.390 140.930 41.670 ;
        RECT 140.720 32.390 140.950 41.390 ;
        RECT 141.855 32.370 142.380 41.395 ;
        RECT 143.255 41.390 143.430 41.670 ;
        RECT 143.580 41.595 144.540 41.825 ;
        RECT 145.030 41.420 145.555 43.720 ;
        RECT 144.630 41.390 145.555 41.420 ;
        RECT 143.255 32.395 143.530 41.390 ;
        RECT 143.300 32.390 143.530 32.395 ;
        RECT 144.590 32.390 145.555 41.390 ;
        RECT 144.630 32.370 145.555 32.390 ;
        RECT 146.880 41.420 147.405 43.720 ;
        RECT 147.880 41.825 148.730 43.245 ;
        RECT 147.880 41.595 148.840 41.825 ;
        RECT 148.980 41.670 156.755 41.845 ;
        RECT 157.005 41.825 157.855 43.245 ;
        RECT 146.880 32.370 148.730 41.420 ;
        RECT 148.980 41.390 149.155 41.670 ;
        RECT 148.890 32.390 149.155 41.390 ;
        RECT 148.980 32.370 149.155 32.390 ;
        RECT 150.030 32.370 150.555 41.395 ;
        RECT 151.505 41.390 151.680 41.670 ;
        RECT 151.470 32.390 151.700 41.390 ;
        RECT 152.605 32.370 153.130 41.395 ;
        RECT 154.080 41.390 154.255 41.670 ;
        RECT 154.050 32.390 154.280 41.390 ;
        RECT 155.180 32.370 155.705 41.395 ;
        RECT 156.580 41.390 156.755 41.670 ;
        RECT 156.910 41.595 157.870 41.825 ;
        RECT 158.355 41.420 158.880 43.720 ;
        RECT 157.955 41.390 158.880 41.420 ;
        RECT 156.580 32.395 156.860 41.390 ;
        RECT 156.630 32.390 156.860 32.395 ;
        RECT 157.920 32.390 158.880 41.390 ;
        RECT 157.955 32.370 158.880 32.390 ;
        RECT 160.205 41.420 160.730 43.720 ;
        RECT 161.205 41.825 162.055 43.245 ;
        RECT 161.205 41.595 162.165 41.825 ;
        RECT 162.305 41.670 170.080 41.845 ;
        RECT 170.330 41.825 171.180 43.245 ;
        RECT 160.205 32.370 162.055 41.420 ;
        RECT 162.305 41.390 162.480 41.670 ;
        RECT 162.215 32.390 162.480 41.390 ;
        RECT 162.305 32.370 162.480 32.390 ;
        RECT 163.355 32.370 163.880 41.395 ;
        RECT 164.830 41.390 165.005 41.670 ;
        RECT 164.795 32.390 165.025 41.390 ;
        RECT 165.930 32.370 166.455 41.395 ;
        RECT 167.405 41.390 167.580 41.670 ;
        RECT 167.375 32.390 167.605 41.390 ;
        RECT 168.505 32.370 169.030 41.395 ;
        RECT 169.905 41.390 170.080 41.670 ;
        RECT 170.235 41.595 171.195 41.825 ;
        RECT 171.680 41.420 172.205 43.720 ;
        RECT 171.280 41.390 172.205 41.420 ;
        RECT 169.905 32.395 170.185 41.390 ;
        RECT 169.955 32.390 170.185 32.395 ;
        RECT 171.245 32.390 172.205 41.390 ;
        RECT 171.280 32.370 172.205 32.390 ;
        RECT 28.905 30.070 29.630 32.370 ;
        RECT 34.395 32.145 35.355 32.185 ;
        RECT 35.685 32.145 36.645 32.185 ;
        RECT 36.975 32.145 37.935 32.185 ;
        RECT 38.265 32.145 39.225 32.185 ;
        RECT 39.555 32.145 40.515 32.185 ;
        RECT 40.845 32.145 41.805 32.185 ;
        RECT 34.395 31.955 41.805 32.145 ;
        RECT 47.720 32.145 48.680 32.185 ;
        RECT 49.010 32.145 49.970 32.185 ;
        RECT 50.300 32.145 51.260 32.185 ;
        RECT 51.590 32.145 52.550 32.185 ;
        RECT 52.880 32.145 53.840 32.185 ;
        RECT 54.170 32.145 55.130 32.185 ;
        RECT 47.720 31.955 55.130 32.145 ;
        RECT 61.045 32.145 62.005 32.185 ;
        RECT 62.335 32.145 63.295 32.185 ;
        RECT 63.625 32.145 64.585 32.185 ;
        RECT 64.915 32.145 65.875 32.185 ;
        RECT 71.795 32.145 72.755 32.185 ;
        RECT 73.085 32.145 74.045 32.185 ;
        RECT 74.375 32.145 75.335 32.185 ;
        RECT 75.665 32.145 76.625 32.185 ;
        RECT 76.955 32.145 77.915 32.185 ;
        RECT 78.245 32.145 79.205 32.185 ;
        RECT 61.045 31.955 65.905 32.145 ;
        RECT 71.795 31.955 79.205 32.145 ;
        RECT 85.120 32.145 86.080 32.185 ;
        RECT 86.410 32.145 87.370 32.185 ;
        RECT 87.700 32.145 88.660 32.185 ;
        RECT 88.990 32.145 89.950 32.185 ;
        RECT 90.280 32.145 91.240 32.185 ;
        RECT 91.570 32.145 92.530 32.185 ;
        RECT 85.120 31.955 92.530 32.145 ;
        RECT 98.445 32.145 99.405 32.185 ;
        RECT 99.735 32.145 100.695 32.185 ;
        RECT 101.025 32.145 101.985 32.185 ;
        RECT 102.315 32.145 103.275 32.185 ;
        RECT 103.605 32.145 104.565 32.185 ;
        RECT 104.895 32.145 105.855 32.185 ;
        RECT 98.445 31.955 105.855 32.145 ;
        RECT 111.770 32.145 112.730 32.185 ;
        RECT 113.060 32.145 114.020 32.185 ;
        RECT 114.350 32.145 115.310 32.185 ;
        RECT 115.640 32.145 116.600 32.185 ;
        RECT 116.930 32.145 117.890 32.185 ;
        RECT 118.220 32.145 119.180 32.185 ;
        RECT 111.770 31.955 119.180 32.145 ;
        RECT 125.095 32.145 126.055 32.185 ;
        RECT 126.385 32.145 127.345 32.185 ;
        RECT 127.675 32.145 128.635 32.185 ;
        RECT 128.965 32.145 129.925 32.185 ;
        RECT 130.255 32.145 131.215 32.185 ;
        RECT 131.545 32.145 132.505 32.185 ;
        RECT 125.095 31.955 132.505 32.145 ;
        RECT 138.420 32.145 139.380 32.185 ;
        RECT 139.710 32.145 140.670 32.185 ;
        RECT 141.000 32.145 141.960 32.185 ;
        RECT 142.290 32.145 143.250 32.185 ;
        RECT 138.420 31.955 143.280 32.145 ;
        RECT 34.405 31.470 41.805 31.955 ;
        RECT 47.730 31.470 55.130 31.955 ;
        RECT 61.055 31.470 65.905 31.955 ;
        RECT 71.805 31.470 79.205 31.955 ;
        RECT 85.130 31.470 92.530 31.955 ;
        RECT 98.455 31.470 105.855 31.955 ;
        RECT 111.780 31.470 119.180 31.955 ;
        RECT 125.105 31.470 132.505 31.955 ;
        RECT 138.430 31.470 143.280 31.955 ;
        RECT 31.555 30.920 41.805 31.470 ;
        RECT 44.880 30.920 55.130 31.470 ;
        RECT 58.205 30.920 65.905 31.470 ;
        RECT 68.955 30.920 79.205 31.470 ;
        RECT 82.280 30.920 92.530 31.470 ;
        RECT 95.605 30.920 105.855 31.470 ;
        RECT 108.930 30.920 119.180 31.470 ;
        RECT 122.255 30.920 132.505 31.470 ;
        RECT 135.580 30.920 143.280 31.470 ;
        RECT 34.405 30.435 41.805 30.920 ;
        RECT 47.730 30.435 55.130 30.920 ;
        RECT 61.055 30.435 65.905 30.920 ;
        RECT 71.805 30.435 79.205 30.920 ;
        RECT 85.130 30.435 92.530 30.920 ;
        RECT 98.455 30.435 105.855 30.920 ;
        RECT 111.780 30.435 119.180 30.920 ;
        RECT 125.105 30.435 132.505 30.920 ;
        RECT 138.430 30.435 143.280 30.920 ;
        RECT 34.395 30.245 41.805 30.435 ;
        RECT 34.395 30.205 35.355 30.245 ;
        RECT 35.685 30.205 36.645 30.245 ;
        RECT 36.975 30.205 37.935 30.245 ;
        RECT 38.265 30.205 39.225 30.245 ;
        RECT 39.555 30.205 40.515 30.245 ;
        RECT 40.845 30.205 41.805 30.245 ;
        RECT 47.720 30.245 55.130 30.435 ;
        RECT 47.720 30.205 48.680 30.245 ;
        RECT 49.010 30.205 49.970 30.245 ;
        RECT 50.300 30.205 51.260 30.245 ;
        RECT 51.590 30.205 52.550 30.245 ;
        RECT 52.880 30.205 53.840 30.245 ;
        RECT 54.170 30.205 55.130 30.245 ;
        RECT 61.045 30.245 65.905 30.435 ;
        RECT 71.795 30.245 79.205 30.435 ;
        RECT 61.045 30.205 62.005 30.245 ;
        RECT 62.335 30.205 63.295 30.245 ;
        RECT 63.625 30.205 64.585 30.245 ;
        RECT 64.915 30.205 65.875 30.245 ;
        RECT 71.795 30.205 72.755 30.245 ;
        RECT 73.085 30.205 74.045 30.245 ;
        RECT 74.375 30.205 75.335 30.245 ;
        RECT 75.665 30.205 76.625 30.245 ;
        RECT 76.955 30.205 77.915 30.245 ;
        RECT 78.245 30.205 79.205 30.245 ;
        RECT 85.120 30.245 92.530 30.435 ;
        RECT 85.120 30.205 86.080 30.245 ;
        RECT 86.410 30.205 87.370 30.245 ;
        RECT 87.700 30.205 88.660 30.245 ;
        RECT 88.990 30.205 89.950 30.245 ;
        RECT 90.280 30.205 91.240 30.245 ;
        RECT 91.570 30.205 92.530 30.245 ;
        RECT 98.445 30.245 105.855 30.435 ;
        RECT 98.445 30.205 99.405 30.245 ;
        RECT 99.735 30.205 100.695 30.245 ;
        RECT 101.025 30.205 101.985 30.245 ;
        RECT 102.315 30.205 103.275 30.245 ;
        RECT 103.605 30.205 104.565 30.245 ;
        RECT 104.895 30.205 105.855 30.245 ;
        RECT 111.770 30.245 119.180 30.435 ;
        RECT 111.770 30.205 112.730 30.245 ;
        RECT 113.060 30.205 114.020 30.245 ;
        RECT 114.350 30.205 115.310 30.245 ;
        RECT 115.640 30.205 116.600 30.245 ;
        RECT 116.930 30.205 117.890 30.245 ;
        RECT 118.220 30.205 119.180 30.245 ;
        RECT 125.095 30.245 132.505 30.435 ;
        RECT 125.095 30.205 126.055 30.245 ;
        RECT 126.385 30.205 127.345 30.245 ;
        RECT 127.675 30.205 128.635 30.245 ;
        RECT 128.965 30.205 129.925 30.245 ;
        RECT 130.255 30.205 131.215 30.245 ;
        RECT 131.545 30.205 132.505 30.245 ;
        RECT 138.420 30.245 143.280 30.435 ;
        RECT 138.420 30.205 139.380 30.245 ;
        RECT 139.710 30.205 140.670 30.245 ;
        RECT 141.000 30.205 141.960 30.245 ;
        RECT 142.290 30.205 143.250 30.245 ;
        RECT 21.355 30.045 22.280 30.070 ;
        RECT 21.355 30.000 22.305 30.045 ;
        RECT 18.225 27.100 22.305 30.000 ;
        RECT 21.355 27.045 22.305 27.100 ;
        RECT 23.365 27.045 23.630 30.045 ;
        RECT 24.530 27.045 24.980 30.045 ;
        RECT 25.945 27.045 26.175 30.045 ;
        RECT 27.130 27.045 27.580 30.045 ;
        RECT 28.480 27.045 28.755 30.045 ;
        RECT 28.905 27.095 30.780 30.070 ;
        RECT 29.815 27.045 30.045 27.095 ;
        RECT 21.355 27.020 22.280 27.045 ;
        RECT 21.355 24.775 21.880 27.020 ;
        RECT 22.355 26.655 23.315 26.885 ;
        RECT 23.455 26.770 23.630 27.045 ;
        RECT 25.980 26.770 26.155 27.045 ;
        RECT 28.480 26.770 28.655 27.045 ;
        RECT 22.355 25.245 23.205 26.655 ;
        RECT 23.455 26.595 28.655 26.770 ;
        RECT 28.805 26.655 29.765 26.885 ;
        RECT 28.855 25.245 29.705 26.655 ;
        RECT 20.500 24.770 22.100 24.775 ;
        RECT 30.255 24.770 30.780 27.095 ;
        RECT 32.105 30.045 33.030 30.070 ;
        RECT 43.180 30.045 44.105 30.070 ;
        RECT 32.105 27.045 33.055 30.045 ;
        RECT 34.115 27.045 34.380 30.045 ;
        RECT 35.280 27.045 35.730 30.045 ;
        RECT 36.695 27.045 36.925 30.045 ;
        RECT 37.880 27.045 38.330 30.045 ;
        RECT 39.275 27.045 39.505 30.045 ;
        RECT 40.455 27.045 40.905 30.045 ;
        RECT 41.805 27.045 42.085 30.045 ;
        RECT 43.145 27.045 44.105 30.045 ;
        RECT 32.105 27.020 33.030 27.045 ;
        RECT 32.105 24.770 32.630 27.020 ;
        RECT 33.105 26.655 34.065 26.885 ;
        RECT 34.205 26.770 34.380 27.045 ;
        RECT 36.730 26.770 36.905 27.045 ;
        RECT 39.305 26.770 39.480 27.045 ;
        RECT 41.805 26.770 41.980 27.045 ;
        RECT 43.180 27.020 44.105 27.045 ;
        RECT 33.105 25.245 33.955 26.655 ;
        RECT 34.205 26.595 41.980 26.770 ;
        RECT 42.135 26.655 43.095 26.885 ;
        RECT 42.230 25.245 43.080 26.655 ;
        RECT 43.580 24.770 44.105 27.020 ;
        RECT 45.430 30.045 46.355 30.070 ;
        RECT 56.505 30.045 57.430 30.070 ;
        RECT 45.430 27.045 46.380 30.045 ;
        RECT 47.440 27.045 47.705 30.045 ;
        RECT 48.605 27.045 49.055 30.045 ;
        RECT 50.020 27.045 50.250 30.045 ;
        RECT 51.205 27.045 51.655 30.045 ;
        RECT 52.600 27.045 52.830 30.045 ;
        RECT 53.780 27.045 54.230 30.045 ;
        RECT 55.130 27.045 55.410 30.045 ;
        RECT 56.470 27.045 57.430 30.045 ;
        RECT 45.430 27.020 46.355 27.045 ;
        RECT 45.430 24.770 45.955 27.020 ;
        RECT 46.430 26.655 47.390 26.885 ;
        RECT 47.530 26.770 47.705 27.045 ;
        RECT 50.055 26.770 50.230 27.045 ;
        RECT 52.630 26.770 52.805 27.045 ;
        RECT 55.130 26.770 55.305 27.045 ;
        RECT 56.505 27.020 57.430 27.045 ;
        RECT 46.430 25.245 47.280 26.655 ;
        RECT 47.530 26.595 55.305 26.770 ;
        RECT 55.460 26.655 56.420 26.885 ;
        RECT 55.555 25.245 56.405 26.655 ;
        RECT 56.905 24.770 57.430 27.020 ;
        RECT 58.755 30.045 59.680 30.070 ;
        RECT 67.255 30.045 68.180 30.070 ;
        RECT 58.755 27.045 59.705 30.045 ;
        RECT 60.765 27.045 61.030 30.045 ;
        RECT 61.930 27.045 62.380 30.045 ;
        RECT 63.345 27.045 63.575 30.045 ;
        RECT 64.530 27.045 64.980 30.045 ;
        RECT 65.880 27.045 66.155 30.045 ;
        RECT 67.215 27.045 68.180 30.045 ;
        RECT 58.755 27.020 59.680 27.045 ;
        RECT 58.755 24.770 59.280 27.020 ;
        RECT 59.755 26.655 60.715 26.885 ;
        RECT 60.855 26.770 61.030 27.045 ;
        RECT 63.380 26.770 63.555 27.045 ;
        RECT 65.880 26.770 66.055 27.045 ;
        RECT 67.255 27.020 68.180 27.045 ;
        RECT 59.755 25.245 60.605 26.655 ;
        RECT 60.855 26.595 66.055 26.770 ;
        RECT 66.205 26.655 67.165 26.885 ;
        RECT 66.255 25.245 67.105 26.655 ;
        RECT 67.655 24.770 68.180 27.020 ;
        RECT 69.505 30.045 70.430 30.070 ;
        RECT 80.580 30.045 81.505 30.070 ;
        RECT 69.505 27.045 70.455 30.045 ;
        RECT 71.515 27.045 71.780 30.045 ;
        RECT 74.095 27.045 74.325 30.045 ;
        RECT 76.675 27.045 76.905 30.045 ;
        RECT 79.205 27.045 79.485 30.045 ;
        RECT 80.545 27.045 81.505 30.045 ;
        RECT 69.505 27.020 70.430 27.045 ;
        RECT 69.505 24.770 70.030 27.020 ;
        RECT 70.505 26.655 71.465 26.885 ;
        RECT 71.605 26.770 71.780 27.045 ;
        RECT 74.130 26.770 74.305 27.045 ;
        RECT 76.705 26.770 76.880 27.045 ;
        RECT 79.205 26.770 79.380 27.045 ;
        RECT 80.580 27.020 81.505 27.045 ;
        RECT 70.505 25.245 71.355 26.655 ;
        RECT 71.605 26.595 79.380 26.770 ;
        RECT 79.535 26.655 80.495 26.885 ;
        RECT 79.630 25.245 80.480 26.655 ;
        RECT 80.980 24.770 81.505 27.020 ;
        RECT 82.830 30.045 83.755 30.070 ;
        RECT 93.905 30.045 94.830 30.070 ;
        RECT 82.830 27.045 83.780 30.045 ;
        RECT 84.840 27.045 85.105 30.045 ;
        RECT 87.420 27.045 87.650 30.045 ;
        RECT 90.000 27.045 90.230 30.045 ;
        RECT 92.530 27.045 92.810 30.045 ;
        RECT 93.870 27.045 94.830 30.045 ;
        RECT 82.830 27.020 83.755 27.045 ;
        RECT 82.830 24.770 83.355 27.020 ;
        RECT 83.830 26.655 84.790 26.885 ;
        RECT 84.930 26.770 85.105 27.045 ;
        RECT 87.455 26.770 87.630 27.045 ;
        RECT 90.030 26.770 90.205 27.045 ;
        RECT 92.530 26.770 92.705 27.045 ;
        RECT 93.905 27.020 94.830 27.045 ;
        RECT 83.830 25.245 84.680 26.655 ;
        RECT 84.930 26.595 92.705 26.770 ;
        RECT 92.860 26.655 93.820 26.885 ;
        RECT 92.955 25.245 93.805 26.655 ;
        RECT 94.305 24.770 94.830 27.020 ;
        RECT 96.155 30.045 97.080 30.070 ;
        RECT 107.230 30.045 108.155 30.070 ;
        RECT 96.155 27.045 97.105 30.045 ;
        RECT 98.165 27.045 98.430 30.045 ;
        RECT 100.745 27.045 100.975 30.045 ;
        RECT 103.325 27.045 103.555 30.045 ;
        RECT 105.855 27.045 106.135 30.045 ;
        RECT 107.195 27.045 108.155 30.045 ;
        RECT 96.155 27.020 97.080 27.045 ;
        RECT 96.155 24.770 96.680 27.020 ;
        RECT 97.155 26.655 98.115 26.885 ;
        RECT 98.255 26.770 98.430 27.045 ;
        RECT 100.780 26.770 100.955 27.045 ;
        RECT 103.355 26.770 103.530 27.045 ;
        RECT 105.855 26.770 106.030 27.045 ;
        RECT 107.230 27.020 108.155 27.045 ;
        RECT 97.155 25.245 98.005 26.655 ;
        RECT 98.255 26.595 106.030 26.770 ;
        RECT 106.185 26.655 107.145 26.885 ;
        RECT 106.280 25.245 107.130 26.655 ;
        RECT 107.630 24.770 108.155 27.020 ;
        RECT 109.480 30.045 110.405 30.070 ;
        RECT 120.555 30.045 121.480 30.070 ;
        RECT 109.480 27.045 110.430 30.045 ;
        RECT 111.490 27.045 111.755 30.045 ;
        RECT 114.070 27.045 114.300 30.045 ;
        RECT 116.650 27.045 116.880 30.045 ;
        RECT 119.180 27.045 119.460 30.045 ;
        RECT 120.520 27.045 121.480 30.045 ;
        RECT 109.480 27.020 110.405 27.045 ;
        RECT 109.480 24.770 110.005 27.020 ;
        RECT 110.480 26.655 111.440 26.885 ;
        RECT 111.580 26.770 111.755 27.045 ;
        RECT 114.105 26.770 114.280 27.045 ;
        RECT 116.680 26.770 116.855 27.045 ;
        RECT 119.180 26.770 119.355 27.045 ;
        RECT 120.555 27.020 121.480 27.045 ;
        RECT 110.480 25.245 111.330 26.655 ;
        RECT 111.580 26.595 119.355 26.770 ;
        RECT 119.510 26.655 120.470 26.885 ;
        RECT 119.605 25.245 120.455 26.655 ;
        RECT 120.955 24.770 121.480 27.020 ;
        RECT 122.805 30.045 123.730 30.070 ;
        RECT 133.880 30.045 134.805 30.070 ;
        RECT 122.805 27.045 123.755 30.045 ;
        RECT 124.815 27.045 125.080 30.045 ;
        RECT 125.980 27.045 126.430 30.045 ;
        RECT 127.395 27.045 127.625 30.045 ;
        RECT 128.580 27.045 129.030 30.045 ;
        RECT 129.975 27.045 130.205 30.045 ;
        RECT 131.155 27.045 131.605 30.045 ;
        RECT 132.505 27.045 132.785 30.045 ;
        RECT 133.845 27.045 134.805 30.045 ;
        RECT 122.805 27.020 123.730 27.045 ;
        RECT 122.805 24.770 123.330 27.020 ;
        RECT 123.805 26.655 124.765 26.885 ;
        RECT 124.905 26.770 125.080 27.045 ;
        RECT 127.430 26.770 127.605 27.045 ;
        RECT 130.005 26.770 130.180 27.045 ;
        RECT 132.505 26.770 132.680 27.045 ;
        RECT 133.880 27.020 134.805 27.045 ;
        RECT 123.805 25.245 124.655 26.655 ;
        RECT 124.905 26.595 132.680 26.770 ;
        RECT 132.835 26.655 133.795 26.885 ;
        RECT 132.930 25.245 133.780 26.655 ;
        RECT 134.280 24.770 134.805 27.020 ;
        RECT 136.130 30.045 137.055 30.070 ;
        RECT 144.630 30.045 145.555 30.070 ;
        RECT 136.130 27.045 137.080 30.045 ;
        RECT 138.140 27.045 138.405 30.045 ;
        RECT 139.305 27.045 139.755 30.045 ;
        RECT 140.720 27.045 140.950 30.045 ;
        RECT 141.905 27.045 142.355 30.045 ;
        RECT 143.255 27.045 143.530 30.045 ;
        RECT 144.590 27.045 145.555 30.045 ;
        RECT 136.130 27.020 137.055 27.045 ;
        RECT 136.130 24.770 136.655 27.020 ;
        RECT 137.130 26.655 138.090 26.885 ;
        RECT 138.230 26.770 138.405 27.045 ;
        RECT 140.755 26.770 140.930 27.045 ;
        RECT 143.255 26.770 143.430 27.045 ;
        RECT 144.630 27.020 145.555 27.045 ;
        RECT 137.130 25.245 137.980 26.655 ;
        RECT 138.230 26.595 143.430 26.770 ;
        RECT 143.580 26.655 144.540 26.885 ;
        RECT 143.630 25.245 144.480 26.655 ;
        RECT 145.030 24.770 145.555 27.020 ;
        RECT 146.880 30.045 147.805 30.070 ;
        RECT 157.955 30.045 158.880 30.070 ;
        RECT 146.880 27.045 147.830 30.045 ;
        RECT 148.890 27.045 149.155 30.045 ;
        RECT 150.055 27.045 150.505 30.045 ;
        RECT 151.470 27.045 151.700 30.045 ;
        RECT 152.655 27.045 153.105 30.045 ;
        RECT 154.050 27.045 154.280 30.045 ;
        RECT 155.230 27.045 155.680 30.045 ;
        RECT 156.580 27.045 156.860 30.045 ;
        RECT 157.920 27.045 158.880 30.045 ;
        RECT 146.880 27.020 147.805 27.045 ;
        RECT 146.880 24.770 147.405 27.020 ;
        RECT 147.880 26.655 148.840 26.885 ;
        RECT 148.980 26.770 149.155 27.045 ;
        RECT 151.505 26.770 151.680 27.045 ;
        RECT 154.080 26.770 154.255 27.045 ;
        RECT 156.580 26.770 156.755 27.045 ;
        RECT 157.955 27.020 158.880 27.045 ;
        RECT 147.880 25.245 148.730 26.655 ;
        RECT 148.980 26.595 156.755 26.770 ;
        RECT 156.910 26.655 157.870 26.885 ;
        RECT 157.005 25.245 157.855 26.655 ;
        RECT 158.355 24.770 158.880 27.020 ;
        RECT 160.205 30.045 161.130 30.070 ;
        RECT 171.280 30.045 172.205 30.070 ;
        RECT 160.205 27.045 161.155 30.045 ;
        RECT 162.215 27.045 162.480 30.045 ;
        RECT 163.380 27.045 163.830 30.045 ;
        RECT 164.795 27.045 165.025 30.045 ;
        RECT 165.980 27.045 166.430 30.045 ;
        RECT 167.375 27.045 167.605 30.045 ;
        RECT 168.555 27.045 169.005 30.045 ;
        RECT 169.905 27.045 170.185 30.045 ;
        RECT 171.245 27.045 172.205 30.045 ;
        RECT 160.205 27.020 161.130 27.045 ;
        RECT 160.205 24.770 160.730 27.020 ;
        RECT 161.205 26.655 162.165 26.885 ;
        RECT 162.305 26.770 162.480 27.045 ;
        RECT 164.830 26.770 165.005 27.045 ;
        RECT 167.405 26.770 167.580 27.045 ;
        RECT 169.905 26.770 170.080 27.045 ;
        RECT 171.280 27.020 172.205 27.045 ;
        RECT 161.205 25.245 162.055 26.655 ;
        RECT 162.305 26.595 170.080 26.770 ;
        RECT 170.235 26.655 171.195 26.885 ;
        RECT 170.330 25.245 171.180 26.655 ;
        RECT 171.680 24.770 172.205 27.020 ;
        RECT 20.500 24.025 172.205 24.770 ;
        RECT 21.105 24.020 172.205 24.025 ;
        RECT 58.025 22.710 59.100 23.750 ;
        RECT 44.735 22.675 44.985 22.710 ;
        RECT 45.565 22.675 45.815 22.710 ;
        RECT 46.395 22.675 46.645 22.710 ;
        RECT 47.225 22.675 47.475 22.710 ;
        RECT 48.055 22.675 48.305 22.710 ;
        RECT 48.885 22.675 49.135 22.710 ;
        RECT 49.715 22.675 49.965 22.710 ;
        RECT 50.545 22.675 50.795 22.710 ;
        RECT 51.375 22.675 51.625 22.710 ;
        RECT 52.205 22.675 52.455 22.710 ;
        RECT 53.035 22.675 53.285 22.710 ;
        RECT 53.865 22.675 54.115 22.710 ;
        RECT 54.695 22.675 54.945 22.710 ;
        RECT 55.525 22.675 55.775 22.710 ;
        RECT 56.355 22.675 56.605 22.710 ;
        RECT 57.185 22.675 57.435 22.710 ;
        RECT 58.015 22.675 59.100 22.710 ;
        RECT 59.675 22.675 59.925 22.710 ;
        RECT 60.505 22.675 60.755 22.710 ;
        RECT 61.335 22.675 61.585 22.710 ;
        RECT 62.165 22.675 62.415 22.710 ;
        RECT 62.995 22.675 63.245 22.710 ;
        RECT 63.825 22.675 64.075 22.710 ;
        RECT 64.655 22.675 64.905 22.710 ;
        RECT 65.485 22.675 65.735 22.710 ;
        RECT 66.315 22.675 66.565 22.710 ;
        RECT 67.145 22.675 67.395 22.710 ;
        RECT 67.975 22.675 68.225 22.710 ;
        RECT 68.805 22.675 69.055 22.710 ;
        RECT 69.635 22.675 69.885 22.710 ;
        RECT 70.465 22.675 70.715 22.710 ;
        RECT 71.295 22.675 71.545 22.710 ;
        RECT 72.125 22.675 72.375 22.710 ;
        RECT 72.955 22.675 73.205 22.710 ;
        RECT 73.785 22.675 74.035 22.710 ;
        RECT 74.615 22.675 74.865 22.710 ;
        RECT 75.445 22.675 75.695 22.710 ;
        RECT 76.275 22.675 76.525 22.710 ;
        RECT 77.105 22.675 77.355 22.710 ;
        RECT 77.935 22.675 78.185 22.710 ;
        RECT 78.765 22.675 79.015 22.710 ;
        RECT 79.595 22.675 79.845 22.710 ;
        RECT 80.425 22.675 80.675 22.710 ;
        RECT 81.255 22.675 81.505 22.710 ;
        RECT 82.085 22.675 82.335 22.710 ;
        RECT 82.915 22.675 83.165 22.710 ;
        RECT 83.745 22.675 83.995 22.710 ;
        RECT 84.575 22.675 84.825 22.710 ;
        RECT 85.405 22.675 85.655 22.710 ;
        RECT 86.235 22.675 86.485 22.710 ;
        RECT 87.065 22.675 87.315 22.710 ;
        RECT 87.895 22.675 88.145 22.710 ;
        RECT 88.725 22.675 88.975 22.710 ;
        RECT 89.555 22.675 89.805 22.710 ;
        RECT 90.385 22.675 90.635 22.710 ;
        RECT 91.215 22.675 91.465 22.710 ;
        RECT 92.045 22.675 92.295 22.710 ;
        RECT 92.875 22.675 93.125 22.710 ;
        RECT 93.705 22.675 93.955 22.710 ;
        RECT 94.535 22.675 94.785 22.710 ;
        RECT 95.365 22.675 95.615 22.710 ;
        RECT 96.195 22.675 96.445 22.710 ;
        RECT 97.025 22.675 97.275 22.710 ;
        RECT 97.855 22.675 98.105 22.710 ;
        RECT 98.685 22.675 98.935 22.710 ;
        RECT 99.515 22.675 99.765 22.710 ;
        RECT 100.345 22.675 100.595 22.710 ;
        RECT 101.175 22.675 101.425 22.710 ;
        RECT 102.005 22.675 102.255 22.710 ;
        RECT 102.835 22.675 103.085 22.710 ;
        RECT 103.665 22.675 103.915 22.710 ;
        RECT 104.495 22.675 104.745 22.710 ;
        RECT 105.325 22.675 105.575 22.710 ;
        RECT 106.155 22.675 106.405 22.710 ;
        RECT 106.985 22.675 107.235 22.710 ;
        RECT 107.815 22.675 108.065 22.710 ;
        RECT 108.645 22.675 108.895 22.710 ;
        RECT 109.475 22.675 109.725 22.710 ;
        RECT 110.305 22.675 110.555 22.710 ;
        RECT 111.135 22.675 111.385 22.710 ;
        RECT 111.965 22.675 112.215 22.710 ;
        RECT 112.795 22.675 113.045 22.710 ;
        RECT 113.625 22.675 113.875 22.710 ;
        RECT 114.455 22.675 114.705 22.710 ;
        RECT 115.285 22.675 115.535 22.710 ;
        RECT 116.115 22.675 116.365 22.710 ;
        RECT 116.945 22.675 117.195 22.710 ;
        RECT 117.775 22.675 118.025 22.710 ;
        RECT 118.605 22.675 118.855 22.710 ;
        RECT 119.435 22.675 119.685 22.710 ;
        RECT 120.265 22.675 120.515 22.710 ;
        RECT 121.095 22.675 121.345 22.710 ;
        RECT 121.925 22.675 122.175 22.710 ;
        RECT 122.755 22.675 123.005 22.710 ;
        RECT 123.585 22.675 123.835 22.710 ;
        RECT 124.415 22.675 124.665 22.710 ;
        RECT 125.245 22.675 125.495 22.710 ;
        RECT 44.725 20.650 45.825 22.675 ;
        RECT 46.395 20.650 47.500 22.675 ;
        RECT 48.050 20.650 49.150 22.675 ;
        RECT 49.715 20.650 50.825 22.675 ;
        RECT 51.375 20.650 52.475 22.675 ;
        RECT 53.035 20.650 54.150 22.675 ;
        RECT 54.695 20.650 55.800 22.675 ;
        RECT 56.350 20.650 57.450 22.675 ;
        RECT 58.015 20.650 59.125 22.675 ;
        RECT 59.675 20.650 60.775 22.675 ;
        RECT 61.335 20.650 62.450 22.675 ;
        RECT 62.995 20.650 64.100 22.675 ;
        RECT 64.650 20.650 65.750 22.675 ;
        RECT 66.315 20.650 67.425 22.675 ;
        RECT 67.975 20.650 69.075 22.675 ;
        RECT 69.635 20.650 70.750 22.675 ;
        RECT 71.295 20.650 72.400 22.675 ;
        RECT 72.955 20.650 74.075 22.675 ;
        RECT 74.615 20.650 75.725 22.675 ;
        RECT 76.275 20.650 77.375 22.675 ;
        RECT 77.935 20.650 79.050 22.675 ;
        RECT 79.595 20.650 80.700 22.675 ;
        RECT 81.250 20.650 82.350 22.675 ;
        RECT 82.915 20.650 84.025 22.675 ;
        RECT 84.575 20.650 85.675 22.675 ;
        RECT 86.235 20.650 87.350 22.675 ;
        RECT 87.895 20.650 89.000 22.675 ;
        RECT 89.550 20.650 90.650 22.675 ;
        RECT 91.200 20.650 92.300 22.675 ;
        RECT 92.875 20.650 93.975 22.675 ;
        RECT 94.535 20.650 95.650 22.675 ;
        RECT 96.195 20.650 97.300 22.675 ;
        RECT 97.850 20.650 98.950 22.675 ;
        RECT 99.515 20.650 100.625 22.675 ;
        RECT 101.175 20.650 102.275 22.675 ;
        RECT 102.825 20.650 103.925 22.675 ;
        RECT 104.495 20.650 105.600 22.675 ;
        RECT 106.150 20.650 107.250 22.675 ;
        RECT 107.815 20.650 108.925 22.675 ;
        RECT 109.475 20.650 110.575 22.675 ;
        RECT 111.135 20.650 112.250 22.675 ;
        RECT 112.795 20.650 113.900 22.675 ;
        RECT 114.450 20.650 115.550 22.675 ;
        RECT 116.115 20.650 117.225 22.675 ;
        RECT 117.775 20.650 118.875 22.675 ;
        RECT 119.435 20.650 120.550 22.675 ;
        RECT 121.095 20.650 122.200 22.675 ;
        RECT 122.750 20.650 123.850 22.675 ;
        RECT 124.415 20.650 125.525 22.675 ;
        RECT 125.900 20.650 126.500 23.750 ;
        RECT 126.725 20.650 127.325 23.225 ;
        RECT 127.735 22.675 127.985 22.710 ;
        RECT 128.565 22.675 128.815 22.710 ;
        RECT 129.395 22.675 129.645 22.710 ;
        RECT 130.225 22.675 130.475 22.710 ;
        RECT 131.055 22.675 131.305 22.710 ;
        RECT 131.885 22.675 132.135 22.710 ;
        RECT 132.715 22.675 132.965 22.710 ;
        RECT 133.545 22.675 133.795 22.710 ;
        RECT 134.375 22.675 134.625 22.710 ;
        RECT 135.205 22.675 135.455 22.710 ;
        RECT 136.035 22.675 136.285 22.710 ;
        RECT 136.865 22.675 137.115 22.710 ;
        RECT 137.695 22.675 137.945 22.710 ;
        RECT 138.525 22.675 138.775 22.710 ;
        RECT 139.355 22.675 139.605 22.710 ;
        RECT 140.185 22.675 140.435 22.710 ;
        RECT 141.015 22.675 141.265 22.710 ;
        RECT 141.845 22.675 142.095 22.710 ;
        RECT 142.675 22.675 142.925 22.710 ;
        RECT 143.505 22.675 143.755 22.710 ;
        RECT 144.335 22.675 144.585 22.710 ;
        RECT 145.165 22.675 145.415 22.710 ;
        RECT 145.995 22.675 146.245 22.710 ;
        RECT 146.825 22.675 147.075 22.710 ;
        RECT 147.655 22.675 147.905 22.710 ;
        RECT 148.485 22.675 148.735 22.710 ;
        RECT 149.315 22.675 149.565 22.710 ;
        RECT 150.145 22.675 150.395 22.710 ;
        RECT 150.975 22.675 151.225 22.710 ;
        RECT 151.805 22.675 152.055 22.710 ;
        RECT 152.635 22.675 152.885 22.710 ;
        RECT 153.465 22.675 153.715 22.710 ;
        RECT 154.295 22.675 154.545 22.710 ;
        RECT 155.125 22.675 155.375 22.710 ;
        RECT 155.955 22.675 156.205 22.710 ;
        RECT 156.785 22.675 157.035 22.710 ;
        RECT 127.735 20.650 128.850 22.675 ;
        RECT 129.395 20.650 130.500 22.675 ;
        RECT 131.050 20.650 132.150 22.675 ;
        RECT 132.715 20.650 133.825 22.675 ;
        RECT 134.375 20.650 135.475 22.675 ;
        RECT 136.035 20.650 137.150 22.675 ;
        RECT 137.695 20.650 138.800 22.675 ;
        RECT 139.350 20.650 140.450 22.675 ;
        RECT 141.015 20.650 142.125 22.675 ;
        RECT 142.675 20.650 143.775 22.675 ;
        RECT 144.335 20.650 145.450 22.675 ;
        RECT 145.995 20.650 147.100 22.675 ;
        RECT 147.650 20.650 148.750 22.675 ;
        RECT 149.315 20.650 150.425 22.675 ;
        RECT 150.975 20.650 152.075 22.675 ;
        RECT 152.635 20.650 153.750 22.675 ;
        RECT 154.295 20.650 155.400 22.675 ;
        RECT 155.950 20.650 157.050 22.675 ;
        RECT 44.735 20.605 44.985 20.650 ;
        RECT 45.565 20.605 45.815 20.650 ;
        RECT 46.395 20.605 46.645 20.650 ;
        RECT 47.225 20.605 47.475 20.650 ;
        RECT 48.055 20.605 48.305 20.650 ;
        RECT 48.885 20.605 49.135 20.650 ;
        RECT 49.715 20.605 49.965 20.650 ;
        RECT 50.545 20.605 50.795 20.650 ;
        RECT 51.375 20.605 51.625 20.650 ;
        RECT 52.205 20.605 52.455 20.650 ;
        RECT 53.035 20.605 53.285 20.650 ;
        RECT 53.865 20.605 54.115 20.650 ;
        RECT 54.695 20.605 54.945 20.650 ;
        RECT 55.525 20.605 55.775 20.650 ;
        RECT 56.355 20.605 56.605 20.650 ;
        RECT 57.185 20.605 57.435 20.650 ;
        RECT 58.015 20.605 58.265 20.650 ;
        RECT 58.845 20.605 59.095 20.650 ;
        RECT 59.675 20.605 59.925 20.650 ;
        RECT 60.505 20.605 60.755 20.650 ;
        RECT 61.335 20.605 61.585 20.650 ;
        RECT 62.165 20.605 62.415 20.650 ;
        RECT 62.995 20.605 63.245 20.650 ;
        RECT 63.825 20.605 64.075 20.650 ;
        RECT 64.655 20.605 64.905 20.650 ;
        RECT 65.485 20.605 65.735 20.650 ;
        RECT 66.315 20.605 66.565 20.650 ;
        RECT 67.145 20.605 67.395 20.650 ;
        RECT 67.975 20.605 68.225 20.650 ;
        RECT 68.805 20.605 69.055 20.650 ;
        RECT 69.635 20.605 69.885 20.650 ;
        RECT 70.465 20.605 70.715 20.650 ;
        RECT 71.295 20.605 71.545 20.650 ;
        RECT 72.125 20.605 72.375 20.650 ;
        RECT 72.955 20.605 73.205 20.650 ;
        RECT 73.785 20.605 74.035 20.650 ;
        RECT 74.615 20.605 74.865 20.650 ;
        RECT 75.445 20.605 75.695 20.650 ;
        RECT 76.275 20.605 76.525 20.650 ;
        RECT 77.105 20.605 77.355 20.650 ;
        RECT 77.935 20.605 78.185 20.650 ;
        RECT 78.765 20.605 79.015 20.650 ;
        RECT 79.595 20.605 79.845 20.650 ;
        RECT 80.425 20.605 80.675 20.650 ;
        RECT 81.255 20.605 81.505 20.650 ;
        RECT 82.085 20.605 82.335 20.650 ;
        RECT 82.915 20.605 83.165 20.650 ;
        RECT 83.745 20.605 83.995 20.650 ;
        RECT 84.575 20.605 84.825 20.650 ;
        RECT 85.405 20.605 85.655 20.650 ;
        RECT 86.235 20.605 86.485 20.650 ;
        RECT 87.065 20.605 87.315 20.650 ;
        RECT 87.895 20.605 88.145 20.650 ;
        RECT 88.725 20.605 88.975 20.650 ;
        RECT 89.555 20.605 89.805 20.650 ;
        RECT 90.385 20.605 90.635 20.650 ;
        RECT 91.215 20.605 91.465 20.650 ;
        RECT 92.045 20.605 92.295 20.650 ;
        RECT 92.875 20.605 93.125 20.650 ;
        RECT 93.705 20.605 93.955 20.650 ;
        RECT 94.535 20.605 94.785 20.650 ;
        RECT 95.365 20.605 95.615 20.650 ;
        RECT 96.195 20.605 96.445 20.650 ;
        RECT 97.025 20.605 97.275 20.650 ;
        RECT 97.855 20.605 98.105 20.650 ;
        RECT 98.685 20.605 98.935 20.650 ;
        RECT 99.515 20.605 99.765 20.650 ;
        RECT 100.345 20.605 100.595 20.650 ;
        RECT 101.175 20.605 101.425 20.650 ;
        RECT 102.005 20.605 102.255 20.650 ;
        RECT 102.835 20.605 103.085 20.650 ;
        RECT 103.665 20.605 103.915 20.650 ;
        RECT 104.495 20.605 104.745 20.650 ;
        RECT 105.325 20.605 105.575 20.650 ;
        RECT 106.155 20.605 106.405 20.650 ;
        RECT 106.985 20.605 107.235 20.650 ;
        RECT 107.815 20.605 108.065 20.650 ;
        RECT 108.645 20.605 108.895 20.650 ;
        RECT 109.475 20.605 109.725 20.650 ;
        RECT 110.305 20.605 110.555 20.650 ;
        RECT 111.135 20.605 111.385 20.650 ;
        RECT 111.965 20.605 112.215 20.650 ;
        RECT 112.795 20.605 113.045 20.650 ;
        RECT 113.625 20.605 113.875 20.650 ;
        RECT 114.455 20.605 114.705 20.650 ;
        RECT 115.285 20.605 115.535 20.650 ;
        RECT 116.115 20.605 116.365 20.650 ;
        RECT 116.945 20.605 117.195 20.650 ;
        RECT 117.775 20.605 118.025 20.650 ;
        RECT 118.605 20.605 118.855 20.650 ;
        RECT 119.435 20.605 119.685 20.650 ;
        RECT 120.265 20.605 120.515 20.650 ;
        RECT 121.095 20.605 121.345 20.650 ;
        RECT 121.925 20.605 122.175 20.650 ;
        RECT 122.755 20.605 123.005 20.650 ;
        RECT 123.585 20.605 123.835 20.650 ;
        RECT 124.415 20.605 124.665 20.650 ;
        RECT 125.245 20.605 125.495 20.650 ;
        RECT 126.075 20.605 126.325 20.650 ;
        RECT 126.905 20.605 127.155 20.650 ;
        RECT 127.735 20.605 127.985 20.650 ;
        RECT 128.565 20.605 128.815 20.650 ;
        RECT 129.395 20.605 129.645 20.650 ;
        RECT 130.225 20.605 130.475 20.650 ;
        RECT 131.055 20.605 131.305 20.650 ;
        RECT 131.885 20.605 132.135 20.650 ;
        RECT 132.715 20.605 132.965 20.650 ;
        RECT 133.545 20.605 133.795 20.650 ;
        RECT 134.375 20.605 134.625 20.650 ;
        RECT 135.205 20.605 135.455 20.650 ;
        RECT 136.035 20.605 136.285 20.650 ;
        RECT 136.865 20.605 137.115 20.650 ;
        RECT 137.695 20.605 137.945 20.650 ;
        RECT 138.525 20.605 138.775 20.650 ;
        RECT 139.355 20.605 139.605 20.650 ;
        RECT 140.185 20.605 140.435 20.650 ;
        RECT 141.015 20.605 141.265 20.650 ;
        RECT 141.845 20.605 142.095 20.650 ;
        RECT 142.675 20.605 142.925 20.650 ;
        RECT 143.505 20.605 143.755 20.650 ;
        RECT 144.335 20.605 144.585 20.650 ;
        RECT 145.165 20.605 145.415 20.650 ;
        RECT 145.995 20.605 146.245 20.650 ;
        RECT 146.825 20.605 147.075 20.650 ;
        RECT 147.655 20.605 147.905 20.650 ;
        RECT 148.485 20.605 148.735 20.650 ;
        RECT 149.315 20.605 149.565 20.650 ;
        RECT 150.145 20.605 150.395 20.650 ;
        RECT 150.975 20.605 151.225 20.650 ;
        RECT 151.805 20.605 152.055 20.650 ;
        RECT 152.635 20.605 152.885 20.650 ;
        RECT 153.465 20.605 153.715 20.650 ;
        RECT 154.295 20.605 154.545 20.650 ;
        RECT 155.125 20.605 155.375 20.650 ;
        RECT 155.955 20.605 156.205 20.650 ;
        RECT 156.785 20.605 157.035 20.650 ;
        RECT 42.850 19.350 43.550 19.975 ;
        RECT 43.905 18.675 44.155 18.715 ;
        RECT 44.735 18.675 44.985 18.715 ;
        RECT 45.565 18.675 45.815 18.715 ;
        RECT 46.395 18.675 46.645 18.715 ;
        RECT 47.225 18.675 47.475 18.715 ;
        RECT 48.055 18.675 48.305 18.715 ;
        RECT 48.885 18.675 49.135 18.715 ;
        RECT 49.715 18.675 49.965 18.715 ;
        RECT 50.545 18.675 50.795 18.715 ;
        RECT 51.375 18.675 51.625 18.715 ;
        RECT 52.205 18.675 52.455 18.715 ;
        RECT 53.035 18.675 53.285 18.715 ;
        RECT 53.865 18.675 54.115 18.715 ;
        RECT 54.695 18.675 54.945 18.715 ;
        RECT 55.525 18.675 55.775 18.715 ;
        RECT 56.355 18.675 56.605 18.715 ;
        RECT 57.185 18.675 57.435 18.715 ;
        RECT 58.015 18.675 58.265 18.715 ;
        RECT 58.845 18.675 59.095 18.715 ;
        RECT 59.675 18.675 59.925 18.715 ;
        RECT 60.505 18.675 60.755 18.715 ;
        RECT 61.335 18.675 61.585 18.715 ;
        RECT 62.165 18.675 62.415 18.715 ;
        RECT 62.995 18.675 63.245 18.715 ;
        RECT 63.825 18.675 64.075 18.715 ;
        RECT 64.655 18.675 64.905 18.715 ;
        RECT 65.485 18.675 65.735 18.715 ;
        RECT 66.315 18.675 66.565 18.715 ;
        RECT 67.145 18.675 67.395 18.715 ;
        RECT 67.975 18.675 68.225 18.715 ;
        RECT 68.805 18.675 69.055 18.715 ;
        RECT 69.635 18.675 69.885 18.715 ;
        RECT 70.465 18.675 70.715 18.715 ;
        RECT 71.295 18.675 71.545 18.715 ;
        RECT 72.125 18.675 72.375 18.715 ;
        RECT 72.955 18.675 73.205 18.715 ;
        RECT 73.785 18.675 74.035 18.715 ;
        RECT 74.615 18.675 74.865 18.715 ;
        RECT 75.445 18.675 75.695 18.715 ;
        RECT 76.275 18.675 76.525 18.715 ;
        RECT 77.105 18.675 77.355 18.715 ;
        RECT 77.935 18.675 78.185 18.715 ;
        RECT 78.765 18.675 79.015 18.715 ;
        RECT 79.595 18.675 79.845 18.715 ;
        RECT 80.425 18.675 80.675 18.715 ;
        RECT 81.255 18.675 81.505 18.715 ;
        RECT 82.085 18.675 82.335 18.715 ;
        RECT 82.915 18.675 83.165 18.715 ;
        RECT 83.745 18.675 83.995 18.715 ;
        RECT 84.575 18.675 84.825 18.715 ;
        RECT 85.405 18.675 85.655 18.715 ;
        RECT 86.235 18.675 86.485 18.715 ;
        RECT 87.065 18.675 87.315 18.715 ;
        RECT 87.895 18.675 88.145 18.715 ;
        RECT 88.725 18.675 88.975 18.715 ;
        RECT 89.555 18.675 89.805 18.715 ;
        RECT 90.385 18.675 90.635 18.715 ;
        RECT 91.215 18.675 91.465 18.715 ;
        RECT 92.045 18.675 92.295 18.715 ;
        RECT 92.875 18.675 93.125 18.715 ;
        RECT 93.705 18.675 93.955 18.715 ;
        RECT 94.535 18.675 94.785 18.715 ;
        RECT 95.365 18.675 95.615 18.715 ;
        RECT 96.195 18.675 96.445 18.715 ;
        RECT 97.025 18.675 97.275 18.715 ;
        RECT 97.855 18.675 98.105 18.715 ;
        RECT 98.685 18.675 98.935 18.715 ;
        RECT 99.515 18.675 99.765 18.715 ;
        RECT 100.345 18.675 100.595 18.715 ;
        RECT 101.175 18.675 101.425 18.715 ;
        RECT 102.005 18.675 102.255 18.715 ;
        RECT 102.835 18.675 103.085 18.715 ;
        RECT 103.665 18.675 103.915 18.715 ;
        RECT 104.495 18.675 104.745 18.715 ;
        RECT 105.325 18.675 105.575 18.715 ;
        RECT 106.155 18.675 106.405 18.715 ;
        RECT 106.985 18.675 107.235 18.715 ;
        RECT 107.815 18.675 108.065 18.715 ;
        RECT 108.645 18.675 108.895 18.715 ;
        RECT 109.475 18.675 109.725 18.715 ;
        RECT 110.305 18.675 110.555 18.715 ;
        RECT 111.135 18.675 111.385 18.715 ;
        RECT 111.965 18.675 112.215 18.715 ;
        RECT 112.795 18.675 113.045 18.715 ;
        RECT 113.625 18.675 113.875 18.715 ;
        RECT 114.455 18.675 114.705 18.715 ;
        RECT 115.285 18.675 115.535 18.715 ;
        RECT 116.115 18.675 116.365 18.715 ;
        RECT 116.945 18.675 117.195 18.715 ;
        RECT 117.775 18.675 118.025 18.715 ;
        RECT 118.605 18.675 118.855 18.715 ;
        RECT 119.435 18.675 119.685 18.715 ;
        RECT 120.265 18.675 120.515 18.715 ;
        RECT 121.095 18.675 121.345 18.715 ;
        RECT 121.925 18.675 122.175 18.715 ;
        RECT 122.755 18.675 123.005 18.715 ;
        RECT 123.585 18.675 123.835 18.715 ;
        RECT 124.415 18.675 124.665 18.715 ;
        RECT 125.245 18.675 125.495 18.715 ;
        RECT 126.075 18.675 126.325 18.715 ;
        RECT 126.905 18.675 127.155 18.715 ;
        RECT 127.735 18.675 127.985 18.715 ;
        RECT 128.565 18.675 128.815 18.715 ;
        RECT 129.395 18.675 129.645 18.715 ;
        RECT 130.225 18.675 130.475 18.715 ;
        RECT 131.055 18.675 131.305 18.715 ;
        RECT 131.885 18.675 132.135 18.715 ;
        RECT 132.715 18.675 132.965 18.715 ;
        RECT 133.545 18.675 133.795 18.715 ;
        RECT 134.375 18.675 134.625 18.715 ;
        RECT 135.205 18.675 135.455 18.715 ;
        RECT 136.035 18.675 136.285 18.715 ;
        RECT 136.865 18.675 137.115 18.715 ;
        RECT 137.695 18.675 137.945 18.715 ;
        RECT 138.525 18.675 138.775 18.715 ;
        RECT 139.355 18.675 139.605 18.715 ;
        RECT 140.185 18.675 140.435 18.715 ;
        RECT 141.015 18.675 141.265 18.715 ;
        RECT 141.845 18.675 142.095 18.715 ;
        RECT 142.675 18.675 142.925 18.715 ;
        RECT 143.505 18.675 143.755 18.715 ;
        RECT 144.335 18.675 144.585 18.715 ;
        RECT 145.165 18.675 145.415 18.715 ;
        RECT 145.995 18.675 146.245 18.715 ;
        RECT 146.825 18.675 147.075 18.715 ;
        RECT 147.655 18.675 147.905 18.715 ;
        RECT 148.485 18.675 148.735 18.715 ;
        RECT 149.315 18.675 149.565 18.715 ;
        RECT 150.145 18.675 150.395 18.715 ;
        RECT 150.975 18.675 151.225 18.715 ;
        RECT 151.805 18.675 152.055 18.715 ;
        RECT 152.635 18.675 152.885 18.715 ;
        RECT 153.465 18.675 153.715 18.715 ;
        RECT 154.295 18.675 154.545 18.715 ;
        RECT 155.125 18.675 155.375 18.715 ;
        RECT 155.955 18.675 156.205 18.715 ;
        RECT 156.785 18.675 157.035 18.715 ;
        RECT 157.615 18.675 157.865 18.715 ;
        RECT 43.900 16.650 45.000 18.675 ;
        RECT 45.550 16.650 46.675 18.675 ;
        RECT 47.225 16.650 48.325 18.675 ;
        RECT 48.875 16.650 49.975 18.675 ;
        RECT 50.545 16.650 51.650 18.675 ;
        RECT 52.200 16.650 53.300 18.675 ;
        RECT 53.850 16.650 54.950 18.675 ;
        RECT 55.525 16.650 56.625 18.675 ;
        RECT 57.175 16.650 58.275 18.675 ;
        RECT 58.845 16.650 59.950 18.675 ;
        RECT 60.500 16.650 61.600 18.675 ;
        RECT 62.165 16.650 63.275 18.675 ;
        RECT 63.825 16.650 64.925 18.675 ;
        RECT 65.475 16.650 66.575 18.675 ;
        RECT 67.145 16.650 68.250 18.675 ;
        RECT 68.800 16.650 69.900 18.675 ;
        RECT 70.465 16.650 71.575 18.675 ;
        RECT 72.125 16.650 73.225 18.675 ;
        RECT 43.905 16.610 44.155 16.650 ;
        RECT 44.735 16.610 44.985 16.650 ;
        RECT 45.565 16.610 45.815 16.650 ;
        RECT 46.395 16.610 46.645 16.650 ;
        RECT 47.225 16.610 47.475 16.650 ;
        RECT 48.055 16.610 48.305 16.650 ;
        RECT 48.885 16.610 49.135 16.650 ;
        RECT 49.715 16.610 49.965 16.650 ;
        RECT 50.545 16.610 50.795 16.650 ;
        RECT 51.375 16.610 51.625 16.650 ;
        RECT 52.205 16.610 52.455 16.650 ;
        RECT 53.035 16.610 53.285 16.650 ;
        RECT 53.865 16.610 54.115 16.650 ;
        RECT 54.695 16.610 54.945 16.650 ;
        RECT 55.525 16.610 55.775 16.650 ;
        RECT 56.355 16.610 56.605 16.650 ;
        RECT 57.185 16.610 57.435 16.650 ;
        RECT 58.015 16.610 58.265 16.650 ;
        RECT 58.845 16.610 59.095 16.650 ;
        RECT 59.675 16.610 59.925 16.650 ;
        RECT 60.505 16.610 60.755 16.650 ;
        RECT 61.335 16.610 61.585 16.650 ;
        RECT 62.165 16.610 62.415 16.650 ;
        RECT 62.995 16.610 63.245 16.650 ;
        RECT 63.825 16.610 64.075 16.650 ;
        RECT 64.655 16.610 64.905 16.650 ;
        RECT 65.485 16.610 65.735 16.650 ;
        RECT 66.315 16.610 66.565 16.650 ;
        RECT 67.145 16.610 67.395 16.650 ;
        RECT 67.975 16.610 68.225 16.650 ;
        RECT 68.805 16.610 69.055 16.650 ;
        RECT 69.635 16.610 69.885 16.650 ;
        RECT 70.465 16.610 70.715 16.650 ;
        RECT 71.295 16.610 71.545 16.650 ;
        RECT 72.125 16.610 72.375 16.650 ;
        RECT 72.955 16.610 73.205 16.650 ;
        RECT 73.775 15.750 74.875 18.675 ;
        RECT 75.445 16.650 76.550 18.675 ;
        RECT 77.100 16.650 78.200 18.675 ;
        RECT 78.765 16.650 79.875 18.675 ;
        RECT 80.425 16.650 81.525 18.675 ;
        RECT 82.075 16.650 83.175 18.675 ;
        RECT 83.745 16.650 84.850 18.675 ;
        RECT 85.400 16.650 86.500 18.675 ;
        RECT 87.065 16.650 88.175 18.675 ;
        RECT 88.725 16.650 89.825 18.675 ;
        RECT 90.385 16.650 91.500 18.675 ;
        RECT 92.045 16.650 93.150 18.675 ;
        RECT 93.700 16.650 94.800 18.675 ;
        RECT 95.365 16.650 96.475 18.675 ;
        RECT 97.025 16.650 98.125 18.675 ;
        RECT 98.685 16.650 99.800 18.675 ;
        RECT 100.345 16.650 101.450 18.675 ;
        RECT 102.000 16.650 103.100 18.675 ;
        RECT 103.665 16.650 104.775 18.675 ;
        RECT 105.325 16.650 106.425 18.675 ;
        RECT 106.975 16.650 108.075 18.675 ;
        RECT 108.645 16.650 109.750 18.675 ;
        RECT 110.300 16.650 111.400 18.675 ;
        RECT 111.965 16.650 113.075 18.675 ;
        RECT 113.625 16.650 114.725 18.675 ;
        RECT 115.275 16.650 116.375 18.675 ;
        RECT 116.925 16.650 118.025 18.675 ;
        RECT 118.600 16.650 119.700 18.675 ;
        RECT 120.265 16.650 121.375 18.675 ;
        RECT 121.925 16.650 123.025 18.675 ;
        RECT 123.575 16.650 124.675 18.675 ;
        RECT 125.245 16.650 126.350 18.675 ;
        RECT 126.900 16.650 128.000 18.675 ;
        RECT 128.565 16.650 129.675 18.675 ;
        RECT 130.225 16.650 131.325 18.675 ;
        RECT 131.885 16.650 133.000 18.675 ;
        RECT 133.545 16.650 134.650 18.675 ;
        RECT 135.200 16.650 136.300 18.675 ;
        RECT 136.850 16.650 137.950 18.675 ;
        RECT 138.525 16.650 139.625 18.675 ;
        RECT 140.175 16.650 141.275 18.675 ;
        RECT 141.825 16.650 142.925 18.675 ;
        RECT 143.500 16.650 144.600 18.675 ;
        RECT 145.165 16.650 146.275 18.675 ;
        RECT 146.825 16.650 147.925 18.675 ;
        RECT 148.475 16.650 149.575 18.675 ;
        RECT 150.145 16.650 151.250 18.675 ;
        RECT 151.800 16.650 152.900 18.675 ;
        RECT 153.450 16.650 154.550 18.675 ;
        RECT 155.125 16.650 156.225 18.675 ;
        RECT 156.775 16.650 157.875 18.675 ;
        RECT 75.445 16.610 75.695 16.650 ;
        RECT 76.275 16.610 76.525 16.650 ;
        RECT 77.105 16.610 77.355 16.650 ;
        RECT 77.935 16.610 78.185 16.650 ;
        RECT 78.765 16.610 79.015 16.650 ;
        RECT 79.595 16.610 79.845 16.650 ;
        RECT 80.425 16.610 80.675 16.650 ;
        RECT 81.255 16.610 81.505 16.650 ;
        RECT 82.085 16.610 82.335 16.650 ;
        RECT 82.915 16.610 83.165 16.650 ;
        RECT 83.745 16.610 83.995 16.650 ;
        RECT 84.575 16.610 84.825 16.650 ;
        RECT 85.405 16.610 85.655 16.650 ;
        RECT 86.235 16.610 86.485 16.650 ;
        RECT 87.065 16.610 87.315 16.650 ;
        RECT 87.895 16.610 88.145 16.650 ;
        RECT 88.725 16.610 88.975 16.650 ;
        RECT 89.555 16.610 89.805 16.650 ;
        RECT 90.385 16.610 90.635 16.650 ;
        RECT 91.215 16.610 91.465 16.650 ;
        RECT 92.045 16.610 92.295 16.650 ;
        RECT 92.875 16.610 93.125 16.650 ;
        RECT 93.705 16.610 93.955 16.650 ;
        RECT 94.535 16.610 94.785 16.650 ;
        RECT 95.365 16.610 95.615 16.650 ;
        RECT 96.195 16.610 96.445 16.650 ;
        RECT 97.025 16.610 97.275 16.650 ;
        RECT 97.855 16.610 98.105 16.650 ;
        RECT 98.685 16.610 98.935 16.650 ;
        RECT 99.515 16.610 99.765 16.650 ;
        RECT 100.345 16.610 100.595 16.650 ;
        RECT 101.175 16.610 101.425 16.650 ;
        RECT 102.005 16.610 102.255 16.650 ;
        RECT 102.835 16.610 103.085 16.650 ;
        RECT 103.665 16.610 103.915 16.650 ;
        RECT 104.495 16.610 104.745 16.650 ;
        RECT 105.325 16.610 105.575 16.650 ;
        RECT 106.155 16.610 106.405 16.650 ;
        RECT 106.985 16.610 107.235 16.650 ;
        RECT 107.815 16.610 108.065 16.650 ;
        RECT 108.645 16.610 108.895 16.650 ;
        RECT 109.475 16.610 109.725 16.650 ;
        RECT 110.305 16.610 110.555 16.650 ;
        RECT 111.135 16.610 111.385 16.650 ;
        RECT 111.965 16.610 112.215 16.650 ;
        RECT 112.795 16.610 113.045 16.650 ;
        RECT 113.625 16.610 113.875 16.650 ;
        RECT 114.455 16.610 114.705 16.650 ;
        RECT 115.285 16.610 115.535 16.650 ;
        RECT 116.115 16.610 116.365 16.650 ;
        RECT 116.945 16.610 117.195 16.650 ;
        RECT 117.775 16.610 118.025 16.650 ;
        RECT 118.605 16.610 118.855 16.650 ;
        RECT 119.435 16.610 119.685 16.650 ;
        RECT 120.265 16.610 120.515 16.650 ;
        RECT 121.095 16.610 121.345 16.650 ;
        RECT 121.925 16.610 122.175 16.650 ;
        RECT 122.755 16.610 123.005 16.650 ;
        RECT 123.585 16.610 123.835 16.650 ;
        RECT 124.415 16.610 124.665 16.650 ;
        RECT 125.245 16.610 125.495 16.650 ;
        RECT 126.075 16.610 126.325 16.650 ;
        RECT 126.905 16.610 127.155 16.650 ;
        RECT 127.735 16.610 127.985 16.650 ;
        RECT 128.565 16.610 128.815 16.650 ;
        RECT 129.395 16.610 129.645 16.650 ;
        RECT 130.225 16.610 130.475 16.650 ;
        RECT 131.055 16.610 131.305 16.650 ;
        RECT 131.885 16.610 132.135 16.650 ;
        RECT 132.715 16.610 132.965 16.650 ;
        RECT 133.545 16.610 133.795 16.650 ;
        RECT 134.375 16.610 134.625 16.650 ;
        RECT 135.205 16.610 135.455 16.650 ;
        RECT 136.035 16.610 136.285 16.650 ;
        RECT 136.865 16.610 137.115 16.650 ;
        RECT 137.695 16.610 137.945 16.650 ;
        RECT 138.525 16.610 138.775 16.650 ;
        RECT 139.355 16.610 139.605 16.650 ;
        RECT 140.185 16.610 140.435 16.650 ;
        RECT 141.015 16.610 141.265 16.650 ;
        RECT 141.845 16.610 142.095 16.650 ;
        RECT 142.675 16.610 142.925 16.650 ;
        RECT 143.505 16.610 143.755 16.650 ;
        RECT 144.335 16.610 144.585 16.650 ;
        RECT 145.165 16.610 145.415 16.650 ;
        RECT 145.995 16.610 146.245 16.650 ;
        RECT 146.825 16.610 147.075 16.650 ;
        RECT 147.655 16.610 147.905 16.650 ;
        RECT 148.485 16.610 148.735 16.650 ;
        RECT 149.315 16.610 149.565 16.650 ;
        RECT 150.145 16.610 150.395 16.650 ;
        RECT 150.975 16.610 151.225 16.650 ;
        RECT 151.805 16.610 152.055 16.650 ;
        RECT 152.635 16.610 152.885 16.650 ;
        RECT 153.465 16.610 153.715 16.650 ;
        RECT 154.295 16.610 154.545 16.650 ;
        RECT 155.125 16.610 155.375 16.650 ;
        RECT 155.955 16.610 156.205 16.650 ;
        RECT 156.785 16.610 157.035 16.650 ;
        RECT 157.615 16.610 157.865 16.650 ;
        RECT 73.775 15.350 127.325 15.750 ;
      LAYER met2 ;
        RECT 125.900 46.000 126.500 47.725 ;
        RECT 126.725 45.325 127.325 53.200 ;
        RECT 30.950 43.245 31.925 43.250 ;
        RECT 22.355 42.495 29.705 43.245 ;
        RECT 30.950 42.500 171.180 43.245 ;
        RECT 22.355 25.995 23.205 41.420 ;
        RECT 24.505 32.370 25.030 41.395 ;
        RECT 27.080 32.370 27.605 41.395 ;
        RECT 24.655 31.470 24.880 32.370 ;
        RECT 27.230 31.470 27.455 32.370 ;
        RECT 28.855 31.895 29.705 42.495 ;
        RECT 30.955 42.495 171.180 42.500 ;
        RECT 30.955 31.470 31.380 42.495 ;
        RECT 24.655 30.920 31.380 31.470 ;
        RECT 31.555 30.920 32.105 31.470 ;
        RECT 24.655 30.045 24.880 30.920 ;
        RECT 27.230 30.045 27.455 30.920 ;
        RECT 24.530 27.045 24.980 30.045 ;
        RECT 27.130 27.045 27.580 30.045 ;
        RECT 33.105 25.995 33.955 41.420 ;
        RECT 35.255 32.370 35.780 41.395 ;
        RECT 37.830 32.370 38.355 41.395 ;
        RECT 40.405 32.370 40.930 41.395 ;
        RECT 35.405 31.470 35.630 32.370 ;
        RECT 37.980 31.470 38.205 32.370 ;
        RECT 40.555 31.470 40.780 32.370 ;
        RECT 44.280 31.470 44.705 37.320 ;
        RECT 35.405 30.920 44.705 31.470 ;
        RECT 44.880 30.920 45.430 31.470 ;
        RECT 35.405 30.045 35.630 30.920 ;
        RECT 37.980 30.045 38.205 30.920 ;
        RECT 40.555 30.045 40.780 30.920 ;
        RECT 35.280 27.045 35.730 30.045 ;
        RECT 37.880 27.045 38.330 30.045 ;
        RECT 40.455 27.045 40.905 30.045 ;
        RECT 46.430 25.995 47.280 41.420 ;
        RECT 48.580 32.370 49.105 41.395 ;
        RECT 51.155 32.370 51.680 41.395 ;
        RECT 53.730 32.370 54.255 41.395 ;
        RECT 48.730 31.470 48.955 32.370 ;
        RECT 51.305 31.470 51.530 32.370 ;
        RECT 53.880 31.470 54.105 32.370 ;
        RECT 57.605 31.470 58.030 37.320 ;
        RECT 48.730 30.920 58.755 31.470 ;
        RECT 48.730 30.045 48.955 30.920 ;
        RECT 51.305 30.045 51.530 30.920 ;
        RECT 53.880 30.045 54.105 30.920 ;
        RECT 48.605 27.045 49.055 30.045 ;
        RECT 51.205 27.045 51.655 30.045 ;
        RECT 53.780 27.045 54.230 30.045 ;
        RECT 59.755 25.995 60.605 41.420 ;
        RECT 61.905 32.370 62.430 41.395 ;
        RECT 64.480 32.370 65.005 41.395 ;
        RECT 62.055 31.470 62.280 32.370 ;
        RECT 64.630 31.470 64.855 32.370 ;
        RECT 62.055 30.920 68.755 31.470 ;
        RECT 68.955 30.920 69.505 31.470 ;
        RECT 62.055 30.045 62.280 30.920 ;
        RECT 64.630 30.045 64.855 30.920 ;
        RECT 68.330 30.145 68.755 30.920 ;
        RECT 61.930 27.045 62.380 30.045 ;
        RECT 64.530 27.045 64.980 30.045 ;
        RECT 70.505 25.995 71.355 41.420 ;
        RECT 82.280 30.920 82.830 31.470 ;
        RECT 83.830 25.995 84.680 41.420 ;
        RECT 95.605 30.920 96.155 31.470 ;
        RECT 97.155 25.995 98.005 41.420 ;
        RECT 108.930 30.920 109.480 31.470 ;
        RECT 110.480 25.995 111.330 41.420 ;
        RECT 122.255 30.920 122.805 31.470 ;
        RECT 123.805 25.995 124.655 41.420 ;
        RECT 125.955 32.370 126.480 41.395 ;
        RECT 128.530 32.370 129.055 41.395 ;
        RECT 131.105 32.370 131.630 41.395 ;
        RECT 126.105 31.470 126.330 32.370 ;
        RECT 128.680 31.470 128.905 32.370 ;
        RECT 131.255 31.470 131.480 32.370 ;
        RECT 134.980 31.470 135.405 33.270 ;
        RECT 126.105 30.920 135.405 31.470 ;
        RECT 135.580 30.920 136.130 31.470 ;
        RECT 126.105 30.045 126.330 30.920 ;
        RECT 128.680 30.045 128.905 30.920 ;
        RECT 131.255 30.045 131.480 30.920 ;
        RECT 125.980 27.045 126.430 30.045 ;
        RECT 128.580 27.045 129.030 30.045 ;
        RECT 131.155 27.045 131.605 30.045 ;
        RECT 137.130 25.995 137.980 41.420 ;
        RECT 139.280 32.370 139.805 41.395 ;
        RECT 141.855 32.370 142.380 41.395 ;
        RECT 139.430 31.470 139.655 32.370 ;
        RECT 142.005 31.470 142.230 32.370 ;
        RECT 139.430 30.920 145.630 31.470 ;
        RECT 139.430 30.045 139.655 30.920 ;
        RECT 142.005 30.045 142.230 30.920 ;
        RECT 139.305 27.045 139.755 30.045 ;
        RECT 141.905 27.045 142.355 30.045 ;
        RECT 147.880 25.995 148.730 41.420 ;
        RECT 150.030 32.370 150.555 41.395 ;
        RECT 152.605 32.370 153.130 41.395 ;
        RECT 155.180 32.370 155.705 41.395 ;
        RECT 150.180 31.470 150.405 32.370 ;
        RECT 152.755 31.470 152.980 32.370 ;
        RECT 155.330 31.470 155.555 32.370 ;
        RECT 159.055 31.470 159.480 37.320 ;
        RECT 150.180 30.920 159.480 31.470 ;
        RECT 150.180 30.045 150.405 30.920 ;
        RECT 152.755 30.045 152.980 30.920 ;
        RECT 155.330 30.045 155.555 30.920 ;
        RECT 150.055 27.045 150.505 30.045 ;
        RECT 152.655 27.045 153.105 30.045 ;
        RECT 155.230 27.045 155.680 30.045 ;
        RECT 161.205 25.995 162.055 41.420 ;
        RECT 163.355 32.370 163.880 41.395 ;
        RECT 165.930 32.370 166.455 41.395 ;
        RECT 168.505 32.370 169.030 41.395 ;
        RECT 163.505 31.470 163.730 32.370 ;
        RECT 166.080 31.470 166.305 32.370 ;
        RECT 168.655 31.470 168.880 32.370 ;
        RECT 172.380 31.470 172.805 37.320 ;
        RECT 163.505 30.920 172.805 31.470 ;
        RECT 163.505 30.045 163.730 30.920 ;
        RECT 166.080 30.045 166.305 30.920 ;
        RECT 168.655 30.045 168.880 30.920 ;
        RECT 163.380 27.045 163.830 30.045 ;
        RECT 165.980 27.045 166.430 30.045 ;
        RECT 168.555 27.045 169.005 30.045 ;
        RECT 22.355 25.245 29.705 25.995 ;
        RECT 33.105 25.245 43.080 25.995 ;
        RECT 46.430 25.245 56.405 25.995 ;
        RECT 59.755 25.245 67.105 25.995 ;
        RECT 70.505 25.245 80.480 25.995 ;
        RECT 83.830 25.245 93.805 25.995 ;
        RECT 97.155 25.245 107.130 25.995 ;
        RECT 110.480 25.245 120.455 25.995 ;
        RECT 123.805 25.245 133.780 25.995 ;
        RECT 137.130 25.245 144.480 25.995 ;
        RECT 147.880 25.245 157.855 25.995 ;
        RECT 161.205 25.245 171.180 25.995 ;
        RECT 42.850 19.350 43.550 24.775 ;
        RECT 125.900 20.800 126.500 22.525 ;
        RECT 126.725 15.350 127.325 23.225 ;
      LAYER met3 ;
        RECT 68.500 46.000 126.500 47.725 ;
        RECT 68.500 44.950 69.325 46.000 ;
        RECT 21.100 43.720 69.325 44.950 ;
        RECT 21.100 43.225 69.330 43.720 ;
        RECT 31.505 31.470 31.930 43.225 ;
        RECT 44.280 36.895 58.030 37.320 ;
        RECT 31.505 30.920 32.105 31.470 ;
        RECT 37.925 25.250 42.530 35.555 ;
        RECT 68.905 31.470 69.330 43.225 ;
        RECT 159.055 36.895 172.805 37.320 ;
        RECT 75.280 32.845 135.405 33.270 ;
        RECT 44.830 30.920 45.430 31.470 ;
        RECT 68.905 30.920 69.505 31.470 ;
        RECT 44.830 25.250 45.255 30.920 ;
        RECT 68.330 29.545 68.755 30.570 ;
        RECT 75.280 29.545 75.730 32.845 ;
        RECT 95.555 31.470 95.980 32.845 ;
        RECT 108.880 31.470 109.305 32.845 ;
        RECT 68.330 29.120 75.730 29.545 ;
        RECT 82.230 30.920 82.830 31.470 ;
        RECT 95.555 30.920 96.155 31.470 ;
        RECT 108.880 30.920 109.480 31.470 ;
        RECT 122.205 30.920 122.805 31.470 ;
        RECT 135.530 30.920 136.130 31.470 ;
        RECT 152.655 30.920 159.055 31.470 ;
        RECT 82.230 25.250 82.655 30.920 ;
        RECT 122.205 29.545 122.630 30.920 ;
        RECT 135.530 29.545 135.955 30.920 ;
        RECT 152.655 29.545 153.105 30.920 ;
        RECT 122.205 29.120 153.105 29.545 ;
        RECT 21.100 24.770 82.655 25.250 ;
        RECT 21.100 23.575 82.650 24.770 ;
        RECT 37.925 11.900 42.530 23.575 ;
        RECT 81.800 22.525 82.650 23.575 ;
        RECT 81.800 20.800 126.500 22.525 ;
  END
END tt_um_TinyWhisper
END LIBRARY

