magic
tech sky130A
magscale 1 2
timestamp 1762799305
<< pwell >>
rect -2196 -20973 2196 20973
<< nmos >>
rect -2000 15763 2000 20763
rect -2000 10545 2000 15545
rect -2000 5327 2000 10327
rect -2000 109 2000 5109
rect -2000 -5109 2000 -109
rect -2000 -10327 2000 -5327
rect -2000 -15545 2000 -10545
rect -2000 -20763 2000 -15763
<< ndiff >>
rect -2058 20751 -2000 20763
rect -2058 15775 -2046 20751
rect -2012 15775 -2000 20751
rect -2058 15763 -2000 15775
rect 2000 20751 2058 20763
rect 2000 15775 2012 20751
rect 2046 15775 2058 20751
rect 2000 15763 2058 15775
rect -2058 15533 -2000 15545
rect -2058 10557 -2046 15533
rect -2012 10557 -2000 15533
rect -2058 10545 -2000 10557
rect 2000 15533 2058 15545
rect 2000 10557 2012 15533
rect 2046 10557 2058 15533
rect 2000 10545 2058 10557
rect -2058 10315 -2000 10327
rect -2058 5339 -2046 10315
rect -2012 5339 -2000 10315
rect -2058 5327 -2000 5339
rect 2000 10315 2058 10327
rect 2000 5339 2012 10315
rect 2046 5339 2058 10315
rect 2000 5327 2058 5339
rect -2058 5097 -2000 5109
rect -2058 121 -2046 5097
rect -2012 121 -2000 5097
rect -2058 109 -2000 121
rect 2000 5097 2058 5109
rect 2000 121 2012 5097
rect 2046 121 2058 5097
rect 2000 109 2058 121
rect -2058 -121 -2000 -109
rect -2058 -5097 -2046 -121
rect -2012 -5097 -2000 -121
rect -2058 -5109 -2000 -5097
rect 2000 -121 2058 -109
rect 2000 -5097 2012 -121
rect 2046 -5097 2058 -121
rect 2000 -5109 2058 -5097
rect -2058 -5339 -2000 -5327
rect -2058 -10315 -2046 -5339
rect -2012 -10315 -2000 -5339
rect -2058 -10327 -2000 -10315
rect 2000 -5339 2058 -5327
rect 2000 -10315 2012 -5339
rect 2046 -10315 2058 -5339
rect 2000 -10327 2058 -10315
rect -2058 -10557 -2000 -10545
rect -2058 -15533 -2046 -10557
rect -2012 -15533 -2000 -10557
rect -2058 -15545 -2000 -15533
rect 2000 -10557 2058 -10545
rect 2000 -15533 2012 -10557
rect 2046 -15533 2058 -10557
rect 2000 -15545 2058 -15533
rect -2058 -15775 -2000 -15763
rect -2058 -20751 -2046 -15775
rect -2012 -20751 -2000 -15775
rect -2058 -20763 -2000 -20751
rect 2000 -15775 2058 -15763
rect 2000 -20751 2012 -15775
rect 2046 -20751 2058 -15775
rect 2000 -20763 2058 -20751
<< ndiffc >>
rect -2046 15775 -2012 20751
rect 2012 15775 2046 20751
rect -2046 10557 -2012 15533
rect 2012 10557 2046 15533
rect -2046 5339 -2012 10315
rect 2012 5339 2046 10315
rect -2046 121 -2012 5097
rect 2012 121 2046 5097
rect -2046 -5097 -2012 -121
rect 2012 -5097 2046 -121
rect -2046 -10315 -2012 -5339
rect 2012 -10315 2046 -5339
rect -2046 -15533 -2012 -10557
rect 2012 -15533 2046 -10557
rect -2046 -20751 -2012 -15775
rect 2012 -20751 2046 -15775
<< psubdiff >>
rect -2160 20903 -2064 20937
rect 2064 20903 2160 20937
rect -2160 20841 -2126 20903
rect 2126 20841 2160 20903
rect -2160 -20903 -2126 -20841
rect 2126 -20903 2160 -20841
rect -2160 -20937 -2064 -20903
rect 2064 -20937 2160 -20903
<< psubdiffcont >>
rect -2064 20903 2064 20937
rect -2160 -20841 -2126 20841
rect 2126 -20841 2160 20841
rect -2064 -20937 2064 -20903
<< poly >>
rect -2000 20835 2000 20851
rect -2000 20801 -1984 20835
rect 1984 20801 2000 20835
rect -2000 20763 2000 20801
rect -2000 15725 2000 15763
rect -2000 15691 -1984 15725
rect 1984 15691 2000 15725
rect -2000 15675 2000 15691
rect -2000 15617 2000 15633
rect -2000 15583 -1984 15617
rect 1984 15583 2000 15617
rect -2000 15545 2000 15583
rect -2000 10507 2000 10545
rect -2000 10473 -1984 10507
rect 1984 10473 2000 10507
rect -2000 10457 2000 10473
rect -2000 10399 2000 10415
rect -2000 10365 -1984 10399
rect 1984 10365 2000 10399
rect -2000 10327 2000 10365
rect -2000 5289 2000 5327
rect -2000 5255 -1984 5289
rect 1984 5255 2000 5289
rect -2000 5239 2000 5255
rect -2000 5181 2000 5197
rect -2000 5147 -1984 5181
rect 1984 5147 2000 5181
rect -2000 5109 2000 5147
rect -2000 71 2000 109
rect -2000 37 -1984 71
rect 1984 37 2000 71
rect -2000 21 2000 37
rect -2000 -37 2000 -21
rect -2000 -71 -1984 -37
rect 1984 -71 2000 -37
rect -2000 -109 2000 -71
rect -2000 -5147 2000 -5109
rect -2000 -5181 -1984 -5147
rect 1984 -5181 2000 -5147
rect -2000 -5197 2000 -5181
rect -2000 -5255 2000 -5239
rect -2000 -5289 -1984 -5255
rect 1984 -5289 2000 -5255
rect -2000 -5327 2000 -5289
rect -2000 -10365 2000 -10327
rect -2000 -10399 -1984 -10365
rect 1984 -10399 2000 -10365
rect -2000 -10415 2000 -10399
rect -2000 -10473 2000 -10457
rect -2000 -10507 -1984 -10473
rect 1984 -10507 2000 -10473
rect -2000 -10545 2000 -10507
rect -2000 -15583 2000 -15545
rect -2000 -15617 -1984 -15583
rect 1984 -15617 2000 -15583
rect -2000 -15633 2000 -15617
rect -2000 -15691 2000 -15675
rect -2000 -15725 -1984 -15691
rect 1984 -15725 2000 -15691
rect -2000 -15763 2000 -15725
rect -2000 -20801 2000 -20763
rect -2000 -20835 -1984 -20801
rect 1984 -20835 2000 -20801
rect -2000 -20851 2000 -20835
<< polycont >>
rect -1984 20801 1984 20835
rect -1984 15691 1984 15725
rect -1984 15583 1984 15617
rect -1984 10473 1984 10507
rect -1984 10365 1984 10399
rect -1984 5255 1984 5289
rect -1984 5147 1984 5181
rect -1984 37 1984 71
rect -1984 -71 1984 -37
rect -1984 -5181 1984 -5147
rect -1984 -5289 1984 -5255
rect -1984 -10399 1984 -10365
rect -1984 -10507 1984 -10473
rect -1984 -15617 1984 -15583
rect -1984 -15725 1984 -15691
rect -1984 -20835 1984 -20801
<< locali >>
rect -2160 20903 -2064 20937
rect 2064 20903 2160 20937
rect -2160 20841 -2126 20903
rect 2126 20841 2160 20903
rect -2000 20801 -1984 20835
rect 1984 20801 2000 20835
rect -2046 20751 -2012 20767
rect -2046 15759 -2012 15775
rect 2012 20751 2046 20767
rect 2012 15759 2046 15775
rect -2000 15691 -1984 15725
rect 1984 15691 2000 15725
rect -2000 15583 -1984 15617
rect 1984 15583 2000 15617
rect -2046 15533 -2012 15549
rect -2046 10541 -2012 10557
rect 2012 15533 2046 15549
rect 2012 10541 2046 10557
rect -2000 10473 -1984 10507
rect 1984 10473 2000 10507
rect -2000 10365 -1984 10399
rect 1984 10365 2000 10399
rect -2046 10315 -2012 10331
rect -2046 5323 -2012 5339
rect 2012 10315 2046 10331
rect 2012 5323 2046 5339
rect -2000 5255 -1984 5289
rect 1984 5255 2000 5289
rect -2000 5147 -1984 5181
rect 1984 5147 2000 5181
rect -2046 5097 -2012 5113
rect -2046 105 -2012 121
rect 2012 5097 2046 5113
rect 2012 105 2046 121
rect -2000 37 -1984 71
rect 1984 37 2000 71
rect -2000 -71 -1984 -37
rect 1984 -71 2000 -37
rect -2046 -121 -2012 -105
rect -2046 -5113 -2012 -5097
rect 2012 -121 2046 -105
rect 2012 -5113 2046 -5097
rect -2000 -5181 -1984 -5147
rect 1984 -5181 2000 -5147
rect -2000 -5289 -1984 -5255
rect 1984 -5289 2000 -5255
rect -2046 -5339 -2012 -5323
rect -2046 -10331 -2012 -10315
rect 2012 -5339 2046 -5323
rect 2012 -10331 2046 -10315
rect -2000 -10399 -1984 -10365
rect 1984 -10399 2000 -10365
rect -2000 -10507 -1984 -10473
rect 1984 -10507 2000 -10473
rect -2046 -10557 -2012 -10541
rect -2046 -15549 -2012 -15533
rect 2012 -10557 2046 -10541
rect 2012 -15549 2046 -15533
rect -2000 -15617 -1984 -15583
rect 1984 -15617 2000 -15583
rect -2000 -15725 -1984 -15691
rect 1984 -15725 2000 -15691
rect -2046 -15775 -2012 -15759
rect -2046 -20767 -2012 -20751
rect 2012 -15775 2046 -15759
rect 2012 -20767 2046 -20751
rect -2000 -20835 -1984 -20801
rect 1984 -20835 2000 -20801
rect -2160 -20903 -2126 -20841
rect 2126 -20903 2160 -20841
rect -2160 -20937 -2064 -20903
rect 2064 -20937 2160 -20903
<< viali >>
rect -1984 20801 1984 20835
rect -2046 15775 -2012 20751
rect 2012 15775 2046 20751
rect -1984 15691 1984 15725
rect -1984 15583 1984 15617
rect -2046 10557 -2012 15533
rect 2012 10557 2046 15533
rect -1984 10473 1984 10507
rect -1984 10365 1984 10399
rect -2046 5339 -2012 10315
rect 2012 5339 2046 10315
rect -1984 5255 1984 5289
rect -1984 5147 1984 5181
rect -2046 121 -2012 5097
rect 2012 121 2046 5097
rect -1984 37 1984 71
rect -1984 -71 1984 -37
rect -2046 -5097 -2012 -121
rect 2012 -5097 2046 -121
rect -1984 -5181 1984 -5147
rect -1984 -5289 1984 -5255
rect -2046 -10315 -2012 -5339
rect 2012 -10315 2046 -5339
rect -1984 -10399 1984 -10365
rect -1984 -10507 1984 -10473
rect -2046 -15533 -2012 -10557
rect 2012 -15533 2046 -10557
rect -1984 -15617 1984 -15583
rect -1984 -15725 1984 -15691
rect -2046 -20751 -2012 -15775
rect 2012 -20751 2046 -15775
rect -1984 -20835 1984 -20801
<< metal1 >>
rect -1996 20835 1996 20841
rect -1996 20801 -1984 20835
rect 1984 20801 1996 20835
rect -1996 20795 1996 20801
rect -2052 20751 -2006 20763
rect -2052 15775 -2046 20751
rect -2012 15775 -2006 20751
rect -2052 15763 -2006 15775
rect 2006 20751 2052 20763
rect 2006 15775 2012 20751
rect 2046 15775 2052 20751
rect 2006 15763 2052 15775
rect -1996 15725 1996 15731
rect -1996 15691 -1984 15725
rect 1984 15691 1996 15725
rect -1996 15685 1996 15691
rect -1996 15617 1996 15623
rect -1996 15583 -1984 15617
rect 1984 15583 1996 15617
rect -1996 15577 1996 15583
rect -2052 15533 -2006 15545
rect -2052 10557 -2046 15533
rect -2012 10557 -2006 15533
rect -2052 10545 -2006 10557
rect 2006 15533 2052 15545
rect 2006 10557 2012 15533
rect 2046 10557 2052 15533
rect 2006 10545 2052 10557
rect -1996 10507 1996 10513
rect -1996 10473 -1984 10507
rect 1984 10473 1996 10507
rect -1996 10467 1996 10473
rect -1996 10399 1996 10405
rect -1996 10365 -1984 10399
rect 1984 10365 1996 10399
rect -1996 10359 1996 10365
rect -2052 10315 -2006 10327
rect -2052 5339 -2046 10315
rect -2012 5339 -2006 10315
rect -2052 5327 -2006 5339
rect 2006 10315 2052 10327
rect 2006 5339 2012 10315
rect 2046 5339 2052 10315
rect 2006 5327 2052 5339
rect -1996 5289 1996 5295
rect -1996 5255 -1984 5289
rect 1984 5255 1996 5289
rect -1996 5249 1996 5255
rect -1996 5181 1996 5187
rect -1996 5147 -1984 5181
rect 1984 5147 1996 5181
rect -1996 5141 1996 5147
rect -2052 5097 -2006 5109
rect -2052 121 -2046 5097
rect -2012 121 -2006 5097
rect -2052 109 -2006 121
rect 2006 5097 2052 5109
rect 2006 121 2012 5097
rect 2046 121 2052 5097
rect 2006 109 2052 121
rect -1996 71 1996 77
rect -1996 37 -1984 71
rect 1984 37 1996 71
rect -1996 31 1996 37
rect -1996 -37 1996 -31
rect -1996 -71 -1984 -37
rect 1984 -71 1996 -37
rect -1996 -77 1996 -71
rect -2052 -121 -2006 -109
rect -2052 -5097 -2046 -121
rect -2012 -5097 -2006 -121
rect -2052 -5109 -2006 -5097
rect 2006 -121 2052 -109
rect 2006 -5097 2012 -121
rect 2046 -5097 2052 -121
rect 2006 -5109 2052 -5097
rect -1996 -5147 1996 -5141
rect -1996 -5181 -1984 -5147
rect 1984 -5181 1996 -5147
rect -1996 -5187 1996 -5181
rect -1996 -5255 1996 -5249
rect -1996 -5289 -1984 -5255
rect 1984 -5289 1996 -5255
rect -1996 -5295 1996 -5289
rect -2052 -5339 -2006 -5327
rect -2052 -10315 -2046 -5339
rect -2012 -10315 -2006 -5339
rect -2052 -10327 -2006 -10315
rect 2006 -5339 2052 -5327
rect 2006 -10315 2012 -5339
rect 2046 -10315 2052 -5339
rect 2006 -10327 2052 -10315
rect -1996 -10365 1996 -10359
rect -1996 -10399 -1984 -10365
rect 1984 -10399 1996 -10365
rect -1996 -10405 1996 -10399
rect -1996 -10473 1996 -10467
rect -1996 -10507 -1984 -10473
rect 1984 -10507 1996 -10473
rect -1996 -10513 1996 -10507
rect -2052 -10557 -2006 -10545
rect -2052 -15533 -2046 -10557
rect -2012 -15533 -2006 -10557
rect -2052 -15545 -2006 -15533
rect 2006 -10557 2052 -10545
rect 2006 -15533 2012 -10557
rect 2046 -15533 2052 -10557
rect 2006 -15545 2052 -15533
rect -1996 -15583 1996 -15577
rect -1996 -15617 -1984 -15583
rect 1984 -15617 1996 -15583
rect -1996 -15623 1996 -15617
rect -1996 -15691 1996 -15685
rect -1996 -15725 -1984 -15691
rect 1984 -15725 1996 -15691
rect -1996 -15731 1996 -15725
rect -2052 -15775 -2006 -15763
rect -2052 -20751 -2046 -15775
rect -2012 -20751 -2006 -15775
rect -2052 -20763 -2006 -20751
rect 2006 -15775 2052 -15763
rect 2006 -20751 2012 -15775
rect 2046 -20751 2052 -15775
rect 2006 -20763 2052 -20751
rect -1996 -20801 1996 -20795
rect -1996 -20835 -1984 -20801
rect 1984 -20835 1996 -20801
rect -1996 -20841 1996 -20835
<< labels >>
rlabel psubdiffcont 0 -20920 0 -20920 0 B
port 1 nsew
rlabel ndiffc -2029 -18263 -2029 -18263 0 D0
port 2 nsew
rlabel ndiffc 2029 -18263 2029 -18263 0 S0
port 3 nsew
rlabel polycont 0 -15708 0 -15708 0 G0
port 4 nsew
rlabel ndiffc -2029 -13045 -2029 -13045 0 D1
port 5 nsew
rlabel ndiffc 2029 -13045 2029 -13045 0 S1
port 6 nsew
rlabel polycont 0 -10490 0 -10490 0 G1
port 7 nsew
rlabel ndiffc -2029 -7827 -2029 -7827 0 D2
port 8 nsew
rlabel ndiffc 2029 -7827 2029 -7827 0 S2
port 9 nsew
rlabel polycont 0 -5272 0 -5272 0 G2
port 10 nsew
rlabel ndiffc -2029 -2609 -2029 -2609 0 D3
port 11 nsew
rlabel ndiffc 2029 -2609 2029 -2609 0 S3
port 12 nsew
rlabel polycont 0 -54 0 -54 0 G3
port 13 nsew
rlabel ndiffc -2029 2609 -2029 2609 0 D4
port 14 nsew
rlabel ndiffc 2029 2609 2029 2609 0 S4
port 15 nsew
rlabel polycont 0 5164 0 5164 0 G4
port 16 nsew
rlabel ndiffc -2029 7827 -2029 7827 0 D5
port 17 nsew
rlabel ndiffc 2029 7827 2029 7827 0 S5
port 18 nsew
rlabel polycont 0 10382 0 10382 0 G5
port 19 nsew
rlabel ndiffc -2029 13045 -2029 13045 0 D6
port 20 nsew
rlabel ndiffc 2029 13045 2029 13045 0 S6
port 21 nsew
rlabel polycont 0 15600 0 15600 0 G6
port 22 nsew
rlabel ndiffc -2029 18263 -2029 18263 0 D7
port 23 nsew
rlabel ndiffc 2029 18263 2029 18263 0 S7
port 24 nsew
rlabel polycont 0 20818 0 20818 0 G7
port 25 nsew
<< properties >>
string FIXED_BBOX -2143 -20920 2143 20920
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 25.0 l 20.0 m 8 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
