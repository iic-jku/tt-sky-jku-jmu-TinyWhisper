magic
tech sky130A
magscale 1 2
timestamp 1762641840
<< locali >>
rect -30 8900 23115 8915
rect -30 8085 -15 8900
rect 25 8845 23060 8860
rect 25 8085 40 8845
rect -30 7385 40 8085
rect 23045 8085 23060 8845
rect 23100 8085 23115 8900
rect 23045 7390 23115 8085
rect -30 2335 40 3030
rect -30 1520 -15 2335
rect 25 1575 40 2335
rect 23045 2335 23115 3030
rect 23045 1575 23060 2335
rect 25 1560 23060 1575
rect 23100 1520 23115 2335
rect -30 1505 23115 1520
<< viali >>
rect -15 8860 23100 8900
rect -15 8085 25 8860
rect 23060 8085 23100 8860
rect -15 1560 25 2335
rect 23060 1560 23100 2335
rect -15 1520 23100 1560
<< metal1 >>
rect -30 8900 23115 8915
rect -30 8085 -15 8900
rect 25 8845 23060 8860
rect 25 8085 40 8845
rect 6115 8735 6345 8745
rect 6115 8330 6125 8735
rect 6335 8330 6345 8735
rect 6115 8320 6345 8330
rect -30 8070 40 8085
rect 23045 8085 23060 8845
rect 23100 8085 23115 8900
rect 23045 8070 23115 8085
rect -65 7530 200 7935
rect 2965 7495 3190 7935
rect 16560 7520 16650 7945
rect 16710 7925 16830 7945
rect 16710 7530 16720 7925
rect 16820 7530 16830 7925
rect 23115 7530 23150 7935
rect 16710 7520 16830 7530
rect -65 2485 200 2890
rect 2970 2880 3190 2920
rect 2970 2485 3185 2880
rect 16560 2475 16650 2900
rect 16710 2890 16830 2900
rect 16710 2485 16720 2890
rect 16820 2485 16830 2890
rect 23115 2485 23150 2890
rect 16710 2475 16830 2485
rect -30 2335 40 2350
rect -30 1520 -15 2335
rect 25 1575 40 2335
rect 23045 2335 23115 2350
rect 6115 2090 6345 2100
rect 6115 1685 6125 2090
rect 6335 1685 6345 2090
rect 16745 1685 16830 2090
rect 6115 1675 6345 1685
rect 23045 1575 23060 2335
rect 25 1560 23060 1575
rect 23100 1520 23115 2335
rect -30 1505 23115 1520
<< via1 >>
rect 6125 8330 6335 8735
rect 16720 7530 16820 7925
rect 16720 2485 16820 2890
rect 6125 1685 6335 2090
<< metal2 >>
rect 6115 8735 6345 8745
rect 6115 8330 6125 8735
rect 6335 8330 16830 8735
rect 6115 8320 16830 8330
rect 16710 7925 16830 8320
rect 16710 7530 16720 7925
rect 16820 7530 16830 7925
rect 16710 7520 16830 7530
rect 16710 2890 16830 2900
rect 16710 2485 16720 2890
rect 16820 2485 16830 2890
rect 16710 2100 16830 2485
rect 6115 2090 16830 2100
rect 6115 1685 6125 2090
rect 6335 1685 16830 2090
rect 6115 1675 16830 1685
use resistors_n  resistors_n_0
timestamp 1762641840
transform 1 0 -165 0 1 -5845
box 100 7350 23315 8914
use resistors_p  resistors_p_0
timestamp 1762641840
transform 1 0 0 0 1 0
box -65 7350 23150 8914
<< end >>
