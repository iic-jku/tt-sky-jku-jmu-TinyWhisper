magic
tech sky130A
magscale 1 2
timestamp 1762641840
<< locali >>
rect -130 4680 1755 4695
rect -130 4365 -115 4680
rect 1740 4365 1755 4680
rect -130 4230 1755 4365
rect -130 4065 20 4230
rect -130 2290 -100 4065
rect -60 2290 20 4065
rect -130 2155 20 2290
rect 1600 4065 1755 4230
rect 1600 2290 1680 4065
rect 1720 2290 1755 4065
rect 1600 2155 1755 2290
rect -130 2130 1755 2155
rect -130 2095 20 2130
rect 1600 2095 1755 2130
rect -130 1925 1755 1985
rect -130 1800 20 1925
rect -130 1220 -100 1800
rect -60 1220 20 1800
rect -130 1070 20 1220
rect 1600 1800 1755 1925
rect 1600 1220 1680 1800
rect 1720 1220 1755 1800
rect 1600 1070 1755 1220
rect -130 925 1755 1070
rect -130 620 -115 925
rect 1740 620 1755 925
rect -130 605 1755 620
<< viali >>
rect -115 4365 1740 4680
rect -100 2290 -60 4065
rect 1680 2290 1720 4065
rect -100 1220 -60 1800
rect 1680 1220 1720 1800
rect -115 620 1740 925
<< metal1 >>
rect -130 4680 1755 4695
rect -130 4365 -115 4680
rect 1740 4365 1755 4680
rect -130 4135 1755 4365
rect -130 4065 375 4135
rect -130 2290 -100 4065
rect -60 2290 375 4065
rect -130 2275 375 2290
rect 475 4070 635 4080
rect 475 2285 485 4070
rect 625 2285 635 4070
rect 475 2275 635 2285
rect 730 2275 890 4135
rect 985 4070 1145 4080
rect 985 2285 995 4070
rect 1135 2285 1145 4070
rect 985 2275 1145 2285
rect 1245 4065 1755 4135
rect 1245 2290 1680 4065
rect 1720 2290 1755 4065
rect 1245 2275 1755 2290
rect 330 2195 1300 2230
rect 325 2165 1300 2195
rect -165 1915 1300 2165
rect 325 1885 1300 1915
rect 330 1850 1300 1885
rect -130 1800 380 1810
rect -130 1220 -100 1800
rect -60 1220 380 1800
rect -130 1155 380 1220
rect 475 1800 635 1810
rect 475 1220 485 1800
rect 625 1220 635 1800
rect 475 1210 635 1220
rect 730 1155 890 1810
rect 985 1800 1145 1810
rect 985 1220 995 1800
rect 1135 1220 1145 1800
rect 985 1210 1145 1220
rect 1240 1800 1755 1810
rect 1240 1220 1680 1800
rect 1720 1220 1755 1800
rect 1240 1155 1755 1220
rect -130 925 1755 1155
rect -130 620 -115 925
rect 1740 620 1755 925
rect -130 605 1755 620
<< via1 >>
rect 485 2285 625 4070
rect 995 2285 1135 4070
rect 485 1220 625 1800
rect 995 1220 1135 1800
<< metal2 >>
rect 475 4070 635 4080
rect 475 2285 485 4070
rect 625 2285 635 4070
rect 475 2240 635 2285
rect 985 4070 1145 4080
rect 985 2285 995 4070
rect 1135 2285 1145 4070
rect 985 2240 1145 2285
rect 475 1840 1770 2240
rect 475 1800 635 1840
rect 475 1220 485 1800
rect 625 1220 635 1800
rect 475 1210 635 1220
rect 985 1800 1145 1840
rect 985 1220 995 1800
rect 1135 1220 1145 1800
rect 985 1210 1145 1220
use sky130_fd_pr__nfet_01v8_lvt_XCBGUP__0  sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0
timestamp 1762641840
transform 1 0 811 0 1 1510
box -941 -510 941 510
use sky130_fd_pr__pfet_01v8_lvt_P4JB26__0  sky130_fd_pr__pfet_01v8_lvt_P4JB26_0
timestamp 1762641840
transform 1 0 811 0 1 3179
box -941 -1119 941 1119
<< labels >>
flabel viali 1040 670 1040 670 0 FreeSans 400 0 0 0 VSS
port 10 nsew
flabel viali 965 4610 965 4610 0 FreeSans 400 0 0 0 VDD
port 11 nsew
flabel metal1 -155 2040 -155 2040 0 FreeSans 320 0 0 0 vin
port 12 nsew
flabel metal2 1760 2040 1760 2040 0 FreeSans 320 0 0 0 vout
port 14 nsew
<< end >>
