magic
tech sky130A
magscale 1 2
timestamp 1762641840
<< pwell >>
rect -359 -310 359 310
<< nmos >>
rect -159 -100 -129 100
rect -63 -100 -33 100
rect 33 -100 63 100
rect 129 -100 159 100
<< ndiff >>
rect -221 88 -159 100
rect -221 -88 -209 88
rect -175 -88 -159 88
rect -221 -100 -159 -88
rect -129 88 -63 100
rect -129 -88 -113 88
rect -79 -88 -63 88
rect -129 -100 -63 -88
rect -33 88 33 100
rect -33 -88 -17 88
rect 17 -88 33 88
rect -33 -100 33 -88
rect 63 88 129 100
rect 63 -88 79 88
rect 113 -88 129 88
rect 63 -100 129 -88
rect 159 88 221 100
rect 159 -88 175 88
rect 209 -88 221 88
rect 159 -100 221 -88
<< ndiffc >>
rect -209 -88 -175 88
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect 175 -88 209 88
<< psubdiff >>
rect -323 240 -227 274
rect 227 240 323 274
rect -323 178 -289 240
rect 289 178 323 240
rect -323 -240 -289 -178
rect 289 -240 323 -178
rect -323 -274 -227 -240
rect 227 -274 323 -240
<< psubdiffcont >>
rect -227 240 227 274
rect -323 -178 -289 178
rect 289 -178 323 178
rect -227 -274 227 -240
<< poly >>
rect -80 190 80 210
rect -80 155 -60 190
rect 60 155 80 190
rect -80 135 80 155
rect -159 100 -129 126
rect -63 100 -33 135
rect 33 100 63 135
rect 129 100 159 126
rect -159 -135 -129 -100
rect -63 -126 -33 -100
rect 33 -126 63 -100
rect -235 -155 -129 -135
rect -235 -190 -215 -155
rect -150 -190 -129 -155
rect -235 -210 -129 -190
rect 129 -135 159 -100
rect 129 -155 235 -135
rect 129 -190 150 -155
rect 215 -190 235 -155
rect 129 -210 235 -190
<< polycont >>
rect -60 155 60 190
rect -215 -190 -150 -155
rect 150 -190 215 -155
<< locali >>
rect -360 274 360 310
rect -360 240 -227 274
rect 227 240 360 274
rect -360 178 -289 240
rect -360 -178 -323 178
rect -80 195 80 205
rect -80 150 -65 195
rect 65 150 80 195
rect -80 140 80 150
rect 289 178 360 240
rect -209 88 -175 104
rect -209 -104 -175 -88
rect -113 88 -79 104
rect -113 -104 -79 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 79 88 113 104
rect 79 -104 113 -88
rect 175 88 209 104
rect 175 -104 209 -88
rect -360 -240 -289 -178
rect -235 -150 -130 -140
rect -235 -195 -220 -150
rect -175 -155 -130 -150
rect -150 -190 -130 -155
rect -175 -195 -130 -190
rect -235 -205 -130 -195
rect 130 -150 235 -140
rect 130 -155 175 -150
rect 130 -190 150 -155
rect 130 -195 175 -190
rect 220 -195 235 -150
rect 130 -205 235 -195
rect 323 -178 360 178
rect 289 -240 360 -178
rect -360 -255 -227 -240
rect 227 -255 360 -240
rect -360 -295 -345 -255
rect 345 -295 360 -255
rect -360 -310 360 -295
<< viali >>
rect -65 190 65 195
rect -65 155 -60 190
rect -60 155 60 190
rect 60 155 65 190
rect -65 150 65 155
rect -209 -88 -175 88
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect 175 -88 209 88
rect -220 -155 -175 -150
rect -220 -190 -215 -155
rect -215 -190 -175 -155
rect -220 -195 -175 -190
rect 175 -155 220 -150
rect 175 -190 215 -155
rect 215 -190 220 -155
rect 175 -195 220 -190
rect -345 -274 -227 -255
rect -227 -274 227 -255
rect 227 -274 345 -255
rect -345 -295 345 -274
<< metal1 >>
rect -80 195 80 205
rect -80 150 -65 195
rect 65 150 80 195
rect -80 140 80 150
rect -215 88 -169 100
rect -215 -88 -209 88
rect -175 -88 -169 88
rect -215 -100 -169 -88
rect -119 88 -73 100
rect -119 -88 -113 88
rect -79 -88 -73 88
rect -119 -100 -73 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 73 88 119 100
rect 73 -88 79 88
rect 113 -88 119 88
rect 73 -100 119 -88
rect 169 88 215 100
rect 169 -88 175 88
rect 209 -88 215 88
rect 169 -100 215 -88
rect -235 -150 -160 -140
rect -235 -195 -220 -150
rect -175 -195 -160 -150
rect -235 -205 -160 -195
rect 160 -150 235 -140
rect 160 -195 175 -150
rect 220 -195 235 -150
rect 160 -205 235 -195
rect -360 -255 360 -240
rect -360 -295 -345 -255
rect 345 -295 360 -255
rect -360 -310 360 -295
<< labels >>
rlabel psubdiffcont 0 -257 0 -257 0 B
port 1 nsew
rlabel ndiffc -192 0 -192 0 0 D0
port 2 nsew
rlabel ndiffc -96 0 -96 0 0 S1
port 4 nsew
rlabel ndiffc 0 0 0 0 0 D2
port 6 nsew
rlabel ndiffc 96 0 96 0 0 S3
port 8 nsew
<< properties >>
string FIXED_BBOX -306 -257 306 257
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 0.150 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
