* PEX produced on Mon Nov 10 03:27:00 PM CET 2025 using /foss/tools/sak/iic-pex.sh with m=1 and s=1
* NGSPICE file created from tt_um_TinyWhisper.ext - technology: sky130A

.subckt tt_um_TinyWhisper_pex clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5] ua[6]
+ ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0]
+ uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0]
+ uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0]
+ uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0]
+ uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7] VDPWR VGND
X0 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_63 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_64 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_118 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_117 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X2 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X3 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_131 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_132 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X4 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_126 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_125 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X5 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X6 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=279.66 ps=1.9598k w=3 l=0.15
X7 VDPWR ui_in[4] iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X8 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X9 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X10 VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X11 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X12 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X13 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_11 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_12 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X14 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X15 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X16 VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X17 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=93.22 ps=735.79999 w=1 l=0.15
X18 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X19 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X20 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=29.46 ps=204.67999 w=3 l=0.15
X21 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X22 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_57 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_56 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X23 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_22 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_21 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X24 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_11 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_10 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X25 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X26 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X27 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_65 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_64 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X28 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X29 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X30 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X31 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_10 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_9 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X32 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X33 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X34 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X35 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_34 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_35 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X36 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_20 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_21 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X37 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_63 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_64 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X38 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X39 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X40 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_74 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_75 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X41 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_15 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_14 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X42 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_131 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_132 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X43 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_37 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X44 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_22 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_23 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X45 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_8 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_9 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X46 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X47 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_76 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_77 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X48 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X49 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X50 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_62 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_63 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X51 VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X52 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X53 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_102 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_101 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X54 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_88 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_87 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X55 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_81 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_82 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X56 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=1.27 ps=4.54 w=1 l=0.15
X57 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_90 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_89 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X58 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_76 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_75 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X59 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_130 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_129 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X60 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X61 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=9.82 ps=76.68 w=1 l=0.15
X62 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X63 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X64 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=55.2 ps=372.79999 w=3 l=0.15
X65 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X66 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X67 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X68 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X69 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X70 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_15 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_14 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X71 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X72 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X73 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X74 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X75 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X76 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X77 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_81 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_82 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X78 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X79 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X80 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_26 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_27 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X81 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n ui_in[4] VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X82 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X83 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_52 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_51 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X84 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X85 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=9.82 ps=76.68 w=1 l=0.15
X86 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X87 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X88 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X89 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_40 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_39 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X90 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X91 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X92 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X93 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X94 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=18.4 ps=148.8 w=1 l=0.15
X95 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X96 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X97 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X98 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X99 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X100 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X101 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X102 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X103 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X104 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X105 VGND VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X106 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X107 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X108 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X109 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X110 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X111 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X112 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X113 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X114 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X115 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X116 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X117 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X118 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X119 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X120 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X121 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X122 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X123 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X124 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X125 VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X126 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X127 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X128 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X129 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X130 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X131 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X132 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X133 VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X134 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X135 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X136 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=29.46 ps=204.67999 w=3 l=0.15
X137 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X138 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X139 ui_in[0] VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X140 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X141 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X142 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X143 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=9.82 ps=76.68 w=1 l=0.15
X144 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X145 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X146 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X147 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X148 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X149 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X150 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X151 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X152 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X153 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X154 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X155 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X156 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X157 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X158 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X159 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X160 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X161 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X162 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X163 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X164 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X165 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X166 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X167 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_116 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_115 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X168 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_55 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_56 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X169 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X170 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X171 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_109 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_110 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X172 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X173 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X174 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X175 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_104 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_103 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X176 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X177 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X178 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X179 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_123 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_122 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X180 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_109 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_108 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X181 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=1.27 ps=4.54 w=1 l=0.15
X182 VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X183 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X184 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X185 VGND VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X186 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X187 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X188 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X189 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X190 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X191 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X192 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X193 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X194 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X195 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_55 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_56 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X196 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X197 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_109 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_110 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X198 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_0 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_1 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X199 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X200 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X201 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X202 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_123 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_122 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X203 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_109 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_108 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X204 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X205 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_59 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_60 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X206 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X207 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_74 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_73 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X208 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X209 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_13 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_14 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X210 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_54 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_53 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X211 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X212 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_128 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_127 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X213 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_122 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_121 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X214 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_67 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_68 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X215 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X216 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X217 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X218 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X219 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_118 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_119 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X220 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_59 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_58 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X221 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_113 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_112 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X222 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X223 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X224 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_120 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_121 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X225 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_135 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_134 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X226 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X227 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_128 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_129 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X228 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X229 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X230 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X231 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X232 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X233 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X234 ui_in[2] VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X235 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X236 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X237 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X238 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=9.82 ps=76.68 w=1 l=0.15
X239 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_59 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_60 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X240 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X241 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X242 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_24 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_25 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X243 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_13 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_14 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X244 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X245 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_67 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_68 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X246 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X247 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X248 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X249 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X250 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X251 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_12 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_13 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X252 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X253 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0 ps=0 w=3 l=1
X254 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_59 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_58 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X255 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_38 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_37 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X256 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_24 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_23 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X257 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_113 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_112 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X258 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_92 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_91 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X259 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_31 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_32 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X260 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_78 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_77 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X261 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_18 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X262 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_135 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_134 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X263 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_3 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_4 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X264 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X265 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_26 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_25 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X266 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X267 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_71 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_72 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X268 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_80 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_79 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X269 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_66 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_65 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X270 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_104 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_105 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X271 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_90 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_91 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X272 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_85 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_84 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X273 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_130 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_131 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X274 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X275 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X276 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_71 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_70 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X277 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_92 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_93 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X278 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X279 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_78 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_79 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X280 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_125 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_124 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X281 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_132 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_133 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X282 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X283 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X284 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X285 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X286 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X287 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_123 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_124 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X288 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X289 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X290 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X291 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X292 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X293 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X294 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X295 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X296 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X297 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X298 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X299 VGND VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X300 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X301 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X302 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_31 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_32 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X303 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_18 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X304 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_3 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_4 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X305 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X306 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X307 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_71 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_72 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X308 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X309 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_2 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_1 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X310 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X311 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X312 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_42 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_41 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X313 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X314 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_28 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_27 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X315 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_85 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_84 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X316 VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X317 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_71 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_70 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X318 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_21 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_22 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X319 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_125 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_124 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X320 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X321 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X322 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_30 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_29 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X323 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_16 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_15 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X324 VGND VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X325 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X326 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_54 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_55 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X327 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X328 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X329 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_40 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_41 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X330 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X331 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X332 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_94 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_95 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X333 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_35 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_34 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X334 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_80 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_81 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X335 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X336 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_21 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_20 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X337 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_42 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_43 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X338 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_123 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_124 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X339 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_28 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_29 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X340 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_96 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_97 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X341 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X342 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X343 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_75 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_74 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X344 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_82 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_83 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X345 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_68 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_69 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X346 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X347 VGND VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X348 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X349 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_108 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_107 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X350 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_94 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_93 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X351 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X352 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_101 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_102 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X353 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_87 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_88 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X354 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_96 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_95 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X355 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X356 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_136 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_135 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X357 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X358 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X359 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X360 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_21 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_22 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X361 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X362 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X363 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_35 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_34 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X364 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_21 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_20 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X365 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X366 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_75 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_74 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X367 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X368 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VGND ui_in[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.93 ps=6.62 w=3 l=0.15
X369 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X370 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X371 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X372 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X373 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X374 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_44 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_45 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X375 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_101 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_102 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X376 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X377 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_87 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_88 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X378 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X379 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X380 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_66 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_67 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X381 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_46 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_47 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X382 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_32 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_33 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X383 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X384 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X385 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=29.46 ps=204.67999 w=3 l=0.15
X386 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X387 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_58 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_57 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X388 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X389 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_112 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_111 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X390 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_51 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_52 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X391 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_46 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_45 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X392 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_100 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X393 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X394 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X395 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X396 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X397 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X398 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0 ps=0 w=3 l=1
X399 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X400 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X401 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X402 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X403 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X404 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X405 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X406 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VGND ui_in[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.93 ps=6.62 w=3 l=0.15
X407 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X408 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X409 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=0 ps=0 w=9 l=1
X410 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X411 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X412 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X413 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X414 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X415 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X416 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X417 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X418 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X419 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X420 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X421 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X422 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X423 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X424 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X425 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=29.46 ps=204.67999 w=3 l=0.15
X426 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_51 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_52 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X427 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X428 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X429 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_16 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X430 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X431 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X432 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X433 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_2 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_3 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X434 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X435 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X436 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_4 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_5 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X437 VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X438 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X439 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X440 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_70 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_69 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X441 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X442 VGND VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X443 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X444 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X445 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X446 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X447 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X448 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X449 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X450 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_136 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X451 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X452 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X453 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X454 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X455 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X456 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X457 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X458 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X459 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X460 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X461 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X462 VGND VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X463 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X464 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X465 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X466 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X467 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X468 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X469 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X470 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X471 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X472 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X473 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X474 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X475 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X476 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X477 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X478 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X479 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X480 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X481 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X482 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X483 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X484 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=0 ps=0 w=9 l=1
X485 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_115 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_116 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X486 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X487 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X488 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X489 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X490 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X491 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X492 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X493 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X494 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X495 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X496 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X497 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X498 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X499 VGND VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X500 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X501 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X502 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X503 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X504 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X505 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X506 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X507 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X508 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X509 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X510 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=0 ps=0 w=9 l=1
X511 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X512 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X513 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X514 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X515 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X516 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_115 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_116 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X517 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X518 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X519 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X520 VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X521 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X522 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X523 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X524 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X525 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X526 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X527 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X528 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X529 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X530 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X531 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_134 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_133 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X532 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X533 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_73 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_74 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X534 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X535 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X536 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X537 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_127 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_128 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X538 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X539 VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X540 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_119 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_118 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X541 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X542 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X543 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X544 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X545 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X546 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X547 VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X548 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X549 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X550 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X551 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X552 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X553 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X554 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X555 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_30 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_31 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X556 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_73 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_74 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X557 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_25 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_24 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X558 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_127 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_128 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X559 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X560 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_18 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_19 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X561 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X562 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X563 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X564 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_44 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_43 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X565 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X566 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X567 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_119 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_118 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X568 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_98 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_97 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X569 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_37 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_38 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X570 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_84 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_83 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X571 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X572 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_23 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_24 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X573 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X574 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_91 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_92 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X575 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_77 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_78 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X576 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_86 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_85 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X577 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X578 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_110 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_111 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X579 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X580 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X581 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_105 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_104 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X582 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_91 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_90 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X583 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X584 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_98 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X585 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_131 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_130 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X586 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X587 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X588 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X589 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X590 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X591 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X592 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X593 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X594 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_25 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_24 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X595 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X596 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=0 ps=0 w=9 l=1
X597 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X598 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X599 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_37 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_38 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X600 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X601 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X602 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_23 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_24 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X603 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_91 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_92 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X604 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_77 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_78 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X605 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X606 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X607 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X608 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X609 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X610 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_62 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_61 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X611 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_48 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_47 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X612 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X613 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_2 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X614 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_34 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_33 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X615 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_105 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_104 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X616 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_91 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_90 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X617 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X618 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_41 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_42 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X619 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_27 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_28 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X620 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_131 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_130 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X621 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_50 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_49 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X622 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_35 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X623 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X624 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X625 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X626 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X627 VGND VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X628 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_60 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_61 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X629 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X630 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_114 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_115 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X631 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_55 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_54 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X632 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_100 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_101 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X633 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X634 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_41 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_40 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X635 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_48 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_49 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X636 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X637 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X638 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_116 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_117 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X639 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_95 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_94 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X640 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X641 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_102 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_103 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X642 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X643 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_81 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_80 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X644 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X645 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X646 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X647 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_88 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_89 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X648 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X649 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X650 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X651 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_114 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_113 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X652 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_107 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_108 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X653 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_93 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_94 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X654 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X655 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VGND ui_in[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.93 ps=6.62 w=3 l=0.15
X656 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X657 VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X658 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X659 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X660 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_2 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X661 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X662 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X663 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_41 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_42 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X664 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_27 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_28 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X665 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X666 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X667 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_6 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_7 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X668 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X669 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_55 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_54 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X670 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X671 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X672 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_41 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_40 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X673 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X674 VGND VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X675 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_20 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_19 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X676 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_6 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_5 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X677 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_95 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_94 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X678 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_0 ua[4] VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X679 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X680 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X681 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_81 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_80 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X682 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X683 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_8 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_7 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X684 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_50 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_51 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X685 VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X686 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X687 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_107 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_108 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X688 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_86 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_87 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X689 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_93 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_94 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X690 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_72 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_73 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X691 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_45 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_44 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X692 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X693 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X694 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_126 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_127 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X695 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_52 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_53 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X696 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_38 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_39 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X697 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_67 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_66 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X698 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_106 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_107 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X699 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X700 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X701 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_118 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_117 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X702 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X703 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_57 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_58 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X704 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X705 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X706 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X707 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_111 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_112 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X708 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_126 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_125 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X709 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_120 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_119 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X710 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_106 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_105 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X711 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X712 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X713 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X714 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X715 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X716 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X717 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X718 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X719 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X720 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X721 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_45 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_44 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X722 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X723 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X724 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_10 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_9 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X725 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_67 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_66 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X726 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X727 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X728 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X729 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_12 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_11 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X730 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X731 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_57 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_58 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X732 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X733 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X734 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_37 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X735 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_22 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_23 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X736 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_8 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_9 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X737 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_111 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_112 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X738 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X739 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X740 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_76 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_77 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X741 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X742 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_16 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X743 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_62 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_63 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X744 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_56 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_57 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X745 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_3 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_2 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X746 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X747 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_10 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_11 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X748 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X749 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X750 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_64 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_65 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X751 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X752 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X753 VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X754 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X755 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_90 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_89 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X756 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X757 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X758 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_76 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_75 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X759 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X760 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_130 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_129 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X761 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_69 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_70 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X762 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_64 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_63 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X763 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X764 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X765 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_132 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_131 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X766 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X767 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X768 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X769 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X770 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X771 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X772 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X773 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_136 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X774 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X775 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X776 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X777 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X778 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X779 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X780 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X781 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X782 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X783 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X784 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_16 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X785 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_3 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_2 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X786 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X787 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X788 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X789 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_26 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_27 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X790 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X791 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VGND ui_in[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.93 ps=6.62 w=3 l=0.15
X792 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X793 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_69 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_70 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X794 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X795 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_14 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_15 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X796 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X797 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X798 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X799 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_40 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_39 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X800 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X801 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin ui_in[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X802 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_136 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X803 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X804 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X805 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_82 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_81 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X806 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X807 VGND VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X808 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X809 VGND VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X810 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X811 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X812 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X813 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n ui_in[4] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X814 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X815 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X816 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X817 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X818 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X819 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=3.81 ps=8.54 w=3 l=0.15
X820 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X821 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X822 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X823 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X824 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X825 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X826 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X827 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X828 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X829 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X830 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X831 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X832 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X833 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X834 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X835 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X836 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X837 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X838 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X839 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X840 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X841 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=3.81 ps=8.54 w=3 l=0.15
X842 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X843 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X844 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X845 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X846 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X847 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X848 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X849 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X850 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X851 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_133 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_134 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X852 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X853 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X854 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X855 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X856 VGND VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X857 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X858 VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X859 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X860 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X861 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=1.27 ps=4.54 w=1 l=0.15
X862 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X863 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X864 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X865 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X866 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X867 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X868 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X869 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X870 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X871 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X872 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X873 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X874 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X875 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X876 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X877 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X878 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X879 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_31 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_30 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X880 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_133 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_134 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X881 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X882 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X883 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X884 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X885 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X886 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X887 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_104 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_103 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X888 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_43 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_44 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X889 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X890 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X891 VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X892 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_97 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_98 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X893 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X894 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_83 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_84 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X895 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X896 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X897 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X898 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X899 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X900 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_111 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_110 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X901 VGND VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X902 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X903 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X904 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_31 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_30 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X905 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X906 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n ui_in[4] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X907 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X908 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X909 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X910 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_0 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_1 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X911 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X912 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X913 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_43 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_44 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X914 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X915 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_97 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_98 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X916 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_83 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_84 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X917 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X918 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X919 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X920 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X921 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X922 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X923 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_54 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_53 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X924 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_111 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_110 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X925 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X926 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_122 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_121 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X927 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_61 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_62 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X928 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_47 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_48 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X929 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X930 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_33 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_34 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X931 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_56 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_55 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X932 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X933 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_110 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_109 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X934 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X935 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X936 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X937 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X938 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X939 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X940 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X941 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_120 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_121 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X942 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_61 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_60 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X943 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X944 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X945 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_115 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_114 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X946 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_128 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_129 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X947 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X948 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_122 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_123 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X949 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_101 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_100 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X950 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_108 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_109 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X951 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X952 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X953 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X954 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X955 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X956 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X957 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_113 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_114 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X958 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X959 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X960 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X961 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X962 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X963 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X964 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X965 VGND ui_in[2] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X966 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_61 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_62 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X967 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_47 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_48 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X968 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_33 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_34 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X969 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X970 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_12 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_13 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X971 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X972 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_7 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_6 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X973 VGND VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X974 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X975 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X976 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_61 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_60 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X977 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=1.27 ps=4.54 w=1 l=0.15
X978 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_26 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_25 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X979 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_115 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_114 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X980 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_101 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_100 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X981 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_80 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_79 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X982 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_19 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_20 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X983 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_66 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_65 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X984 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_60 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_59 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X985 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_5 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_6 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X986 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X987 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_14 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_13 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X988 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X989 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VDPWR ui_in[1] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X990 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_68 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_67 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X991 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X992 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_113 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_114 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X993 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_92 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_93 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X994 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X995 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_78 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_79 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X996 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_51 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_50 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X997 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_58 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_59 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X998 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_87 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_86 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X999 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1000 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1001 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_132 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_133 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1002 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_73 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_72 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1003 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1004 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_112 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_113 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1005 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_127 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_126 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1006 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1007 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1008 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_134 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_135 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1009 ui_in[1] VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0.495 ps=3.33 w=3 l=0.15
X1010 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1011 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1012 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1013 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1014 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_117 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_118 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1015 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1016 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1017 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1018 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1019 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_125 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_126 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1020 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1021 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_7 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_6 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1022 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1023 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1024 VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X1025 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1026 VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X1027 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_19 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_20 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1028 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_5 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_6 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1029 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1030 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n ui_in[4] VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1031 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1032 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1033 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1034 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_51 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_50 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1035 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_30 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_29 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1036 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_16 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_15 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1037 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_87 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_86 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1038 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1039 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X1040 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_73 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_72 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1041 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1042 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1043 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1044 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_9 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_10 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1045 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_127 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_126 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1046 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_32 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_31 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1047 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1048 ui_in[3] VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0.495 ps=3.33 w=3 l=0.15
X1049 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_18 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1050 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1051 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_4 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_3 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1052 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_72 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_71 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1053 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1054 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1055 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_42 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_43 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1056 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1057 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_28 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_29 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1058 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_117 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_118 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1059 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1060 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin ui_in[0] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1061 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_96 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_97 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1062 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_37 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1063 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1064 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_82 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_83 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1065 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_23 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_22 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1066 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_68 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_69 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1067 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_125 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_126 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1068 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_9 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_8 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1069 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1070 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1071 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_77 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_76 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1072 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_63 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_62 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1073 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_84 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_85 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1074 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_70 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_71 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1075 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_124 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_125 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1076 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1077 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_96 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_95 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1078 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1079 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_89 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_90 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1080 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_136 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_135 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1081 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_75 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_76 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1082 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1083 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1084 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_129 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_130 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1085 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1086 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_124 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_123 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1087 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1088 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1089 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_9 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_10 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1090 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1091 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1092 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1093 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1094 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1095 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1096 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1097 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1098 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin ui_in[2] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1099 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1100 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_37 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1101 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1102 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_23 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_22 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1103 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1104 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_9 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_8 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1105 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_77 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_76 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1106 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1107 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1108 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_63 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_62 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1109 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1110 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_22 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_21 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1111 VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X1112 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1113 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1114 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_46 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_47 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1115 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_32 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_33 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1116 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1117 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_89 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_90 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1118 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_75 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_76 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1119 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1120 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_27 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_26 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1121 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_129 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_130 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1122 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_34 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_35 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1123 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1124 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_20 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_21 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1125 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1126 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1127 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_74 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_75 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1128 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1129 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1130 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_46 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_45 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1131 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_100 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1132 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_39 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_40 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1133 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=3.81 ps=8.54 w=3 l=0.15
X1134 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1135 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1136 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_102 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_101 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1137 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_88 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_87 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1138 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1139 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1140 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1141 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1142 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1143 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1144 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1145 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VDPWR ui_in[3] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X1146 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1147 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1148 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1149 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1150 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1151 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_27 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_26 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1152 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1153 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1154 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1155 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1156 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1157 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1158 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1159 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_39 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_40 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1160 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1161 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1162 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_4 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_5 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1163 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1164 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1165 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1166 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1167 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1168 VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X1169 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1170 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1171 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_52 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_51 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1172 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1173 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n ui_in[4] VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1174 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1175 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=1.27 ps=4.54 w=1 l=0.15
X1176 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1177 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1178 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1179 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1180 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X1181 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1182 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin ui_in[1] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1183 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1184 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1185 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1186 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1187 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1188 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1189 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1190 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1191 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1192 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1193 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X1194 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1195 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1196 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1197 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1198 VGND ui_in[4] iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1199 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1200 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1201 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1202 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1203 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1204 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1205 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1206 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1207 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin ui_in[3] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1208 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1209 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1210 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1211 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1212 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1213 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1214 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1215 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1216 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1217 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1218 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1219 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1220 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1221 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1222 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1223 VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X1224 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1225 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin ui_in[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1226 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1227 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1228 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_103 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_104 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1229 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1230 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1231 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1232 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1233 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=3.81 ps=8.54 w=3 l=0.15
X1234 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1235 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1236 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1237 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1238 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1239 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1240 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1241 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1242 VDPWR ui_in[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1243 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1244 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1245 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1246 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1247 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1248 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1249 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1250 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1251 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1252 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_0 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1253 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_103 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_104 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1254 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1255 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_53 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_54 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1256 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_121 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_122 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1257 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1258 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1259 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1260 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_116 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_115 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1261 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1262 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1263 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1264 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1265 VDPWR ui_in[2] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1266 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_121 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_120 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1267 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1268 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_129 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_128 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1269 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1270 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1271 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1272 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=1.27 ps=4.54 w=1 l=0.15
X1273 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1274 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1275 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=1.27 ps=4.54 w=1 l=0.15
X1276 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1277 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_0 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1278 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1279 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1280 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1281 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1282 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1283 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VDPWR ui_in[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X1284 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1285 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1286 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1287 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1288 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1289 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1290 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_53 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_54 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1291 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_121 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_122 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1292 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1293 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_18 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_19 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1294 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X1295 ui_in[0] VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0.495 ps=3.33 w=3 l=0.15
X1296 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1297 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_13 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_12 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1298 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1299 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1300 VGND ui_in[4] iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1301 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1302 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_121 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_120 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1303 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1304 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_86 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_85 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1305 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_25 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_26 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1306 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_129 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_128 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1307 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_79 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_80 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1308 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_65 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_66 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1309 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1310 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_74 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_73 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1311 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1312 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1313 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_128 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_127 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1314 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1315 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1316 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_98 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1317 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1318 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1319 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1320 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1321 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_93 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_92 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1322 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1323 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_79 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_78 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1324 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_118 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_119 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1325 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_133 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_132 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1326 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1327 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1328 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1329 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1330 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1331 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1332 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1333 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1334 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_13 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_12 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1335 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1336 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1337 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1338 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1339 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin ui_in[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1340 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_25 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_26 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1341 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1342 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_79 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_80 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1343 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_65 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_66 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1344 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1345 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1346 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_24 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_25 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1347 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_50 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_49 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1348 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_35 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1349 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_93 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_92 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1350 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_79 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_78 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1351 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1352 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_29 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_30 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1353 VDPWR ui_in[1] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1354 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_133 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_132 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1355 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_38 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_37 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1356 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_15 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_16 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1357 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_24 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_23 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1358 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1359 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_92 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_91 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1360 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_78 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_77 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1361 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1362 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_48 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_49 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1363 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_116 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_117 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1364 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1365 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_102 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_103 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1366 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1367 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1368 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_43 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_42 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1369 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_88 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_89 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1370 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_29 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_28 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1371 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_97 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_96 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1372 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_83 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_82 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1373 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1374 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_104 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_105 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1375 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_69 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_68 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1376 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_90 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_91 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1377 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_130 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_131 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1378 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1379 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1380 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_95 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_96 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1381 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1382 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1383 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_135 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_136 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1384 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X1385 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1386 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1387 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1388 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1389 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1390 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1391 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_29 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_30 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1392 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1393 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_15 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_16 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1394 VDPWR ui_in[3] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1395 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1396 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_0 ua[2] VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1397 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_43 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_42 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1398 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_29 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_28 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1399 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_8 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_7 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1400 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_97 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_96 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1401 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_83 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_82 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1402 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1403 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_2 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_1 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1404 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_69 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_68 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1405 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_42 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_41 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1406 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1407 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_28 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_27 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1408 VGND ui_in[1] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1409 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_52 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_53 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1410 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_38 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_39 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1411 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1412 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_106 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_107 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1413 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_95 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_96 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1414 VDPWR ui_in[4] iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1415 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1416 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_47 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_46 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1417 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1418 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_54 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_55 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1419 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_33 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_32 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1420 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_135 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_136 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1421 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_40 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_41 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1422 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1423 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VDPWR ui_in[2] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X1424 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1425 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_94 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_95 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1426 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_80 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_81 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1427 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1428 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_120 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_119 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1429 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_106 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_105 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1430 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_45 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_46 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1431 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1432 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_100 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1433 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1434 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1435 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1436 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_108 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_107 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1437 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1438 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_94 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_93 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1439 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1440 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1441 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1442 ui_in[2] VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0.495 ps=3.33 w=3 l=0.15
X1443 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1444 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1445 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1446 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1447 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1448 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1449 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1450 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1451 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1452 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1453 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1454 VGND ui_in[4] iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1455 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1456 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_47 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_46 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1457 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1458 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_33 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_32 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1459 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1460 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_12 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_11 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1461 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1462 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1463 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_45 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_46 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1464 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_56 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_57 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1465 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1466 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_10 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_11 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1467 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_100 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1468 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1469 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_64 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_65 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1470 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1471 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1472 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_5 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_4 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1473 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_44 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_45 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1474 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1475 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1476 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1477 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_66 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_67 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1478 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1479 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1480 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1481 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_64 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_63 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1482 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_58 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_57 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1483 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_132 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_131 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1484 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1485 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_112 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_111 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1486 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1487 VGND VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X1488 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1489 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1490 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1491 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1492 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1493 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_5 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_4 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1494 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1495 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1496 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1497 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1498 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1499 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1500 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1501 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1502 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1503 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1504 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_14 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_15 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1505 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X1506 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_16 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1507 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_2 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_3 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1508 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1509 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin ui_in[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1510 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1511 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1512 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1513 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1514 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1515 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_82 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_81 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1516 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1517 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1518 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1519 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n ui_in[4] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1520 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X1521 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_70 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_69 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1522 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1523 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1524 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1525 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1526 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_136 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1527 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1528 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1529 VGND ui_in[3] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1530 VDPWR ui_in[4] iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1531 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1532 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1533 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1534 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1535 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1536 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=3.81 ps=8.54 w=3 l=0.15
X1537 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1538 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1539 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1540 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1541 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1542 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1543 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1544 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1545 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1546 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1547 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1548 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1549 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1550 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1551 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1552 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1553 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1554 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1555 VGND ui_in[4] iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1556 VGND VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X1557 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1558 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1559 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1560 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1561 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1562 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=3.81 ps=8.54 w=3 l=0.15
X1563 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1564 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1565 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1566 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1567 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1568 VGND VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X1569 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1570 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1571 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1572 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1573 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1574 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1575 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1576 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1577 VGND VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X1578 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1579 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1580 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1581 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1582 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1583 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1584 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1585 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1586 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1587 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1588 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1589 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_19 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_18 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1590 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1591 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1592 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1593 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_85 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_86 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1594 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_134 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_133 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1595 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1596 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1597 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1598 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_98 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1599 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1600 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1601 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1602 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X1603 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1604 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1605 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n ui_in[4] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1606 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X1607 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1608 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1609 ui_in[1] VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X1610 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1611 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1612 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1613 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1614 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1615 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1616 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_19 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_18 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1617 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=3.81 ps=8.54 w=3 l=0.15
X1618 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1619 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1620 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1621 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_85 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_86 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1622 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_30 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_31 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1623 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1624 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1625 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1626 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1627 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_56 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_55 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1628 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1629 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1630 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1631 VDPWR ui_in[4] iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1632 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_110 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_109 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1633 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_98 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1634 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_49 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_50 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1635 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_35 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1636 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1637 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_44 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_43 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1638 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1639 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_98 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_97 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1640 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_84 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_83 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1641 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1642 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_122 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_123 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1643 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1644 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_108 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_109 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1645 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_49 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_48 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1646 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_117 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_116 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1647 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_103 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_102 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1648 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1649 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_89 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_88 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1650 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_110 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_111 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1651 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1652 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1653 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1654 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1655 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1656 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=3.81 ps=8.54 w=3 l=0.15
X1657 VGND VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X1658 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1659 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1660 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1661 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1662 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1663 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1664 VGND VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X1665 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1666 VGND ui_in[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1667 VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X1668 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1669 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_49 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_50 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1670 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_35 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1671 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=1.27 ps=4.54 w=1 l=0.15
X1672 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1673 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1674 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1675 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1676 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1677 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_49 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_48 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1678 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_60 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_59 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1679 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_117 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_116 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1680 ua[1] iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_0 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1681 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_14 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_13 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1682 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_103 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_102 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1683 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_89 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_88 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1684 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_68 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_67 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1685 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_62 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_61 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1686 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_7 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_8 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1687 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_48 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_47 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1688 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_34 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_33 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1689 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1690 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1691 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_58 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_59 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1692 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_112 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_113 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1693 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1694 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1695 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_53 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_52 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1696 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_60 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_61 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1697 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_39 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_38 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1698 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_134 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_135 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1699 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1700 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1701 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_107 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_106 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1702 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1703 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_114 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_115 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1704 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_100 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_101 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1705 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1706 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1707 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_119 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_120 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1708 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_105 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_106 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1709 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1710 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_114 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_113 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1711 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1712 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n ui_in[4] VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1713 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1714 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1715 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1716 ua[3] iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_0 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1717 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1718 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1719 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1720 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_7 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_8 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1721 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1722 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_6 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_7 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1723 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1724 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1725 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_53 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_52 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1726 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_32 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_31 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1727 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_39 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_38 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1728 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1729 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X1730 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_18 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1731 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_107 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_106 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1732 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_4 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_3 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1733 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1734 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_72 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_71 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1735 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_11 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_12 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1736 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_20 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_19 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1737 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1738 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_6 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_5 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1739 ui_in[3] VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X1740 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1741 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_119 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_120 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1742 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1743 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1744 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_105 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_106 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1745 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1746 VGND VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X1747 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_84 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_85 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1748 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_57 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_56 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1749 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_70 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_71 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1750 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_11 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_10 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1751 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_50 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_51 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1752 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1753 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_124 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_125 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1754 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_65 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_64 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1755 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_86 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_87 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1756 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_72 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_73 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1757 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_126 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_127 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1758 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1759 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1760 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1761 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1762 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_124 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_123 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1763 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
C0 ua[5] VGND 0.14696f
C1 ua[6] VGND 0.14696f
C2 ua[7] VGND 0.14696f
C3 ena VGND 0.09789f
C4 clk VGND 0.09789f
C5 rst_n VGND 0.09789f
C6 ui_in[5] VGND 0.09789f
C7 ui_in[6] VGND 0.09789f
C8 ui_in[7] VGND 0.09789f
C9 uio_in[0] VGND 0.09789f
C10 uio_in[1] VGND 0.09789f
C11 uio_in[2] VGND 0.09789f
C12 uio_in[3] VGND 0.09789f
C13 uio_in[4] VGND 0.09789f
C14 uio_in[5] VGND 0.09789f
C15 uio_in[6] VGND 0.09789f
C16 uio_in[7] VGND 0.09789f
C17 uo_out[0] VGND 0.09789f
C18 uo_out[1] VGND 0.09789f
C19 uo_out[2] VGND 0.09789f
C20 uo_out[3] VGND 0.09789f
C21 uo_out[4] VGND 0.09789f
C22 uo_out[5] VGND 0.09789f
C23 uo_out[6] VGND 0.09789f
C24 uo_out[7] VGND 0.09789f
C25 uio_out[0] VGND 0.09789f
C26 uio_out[1] VGND 0.09789f
C27 uio_out[2] VGND 0.09789f
C28 uio_out[3] VGND 0.09789f
C29 uio_out[4] VGND 0.09789f
C30 uio_out[5] VGND 0.09789f
C31 uio_out[6] VGND 0.09789f
C32 uio_out[7] VGND 0.09789f
C33 uio_oe[0] VGND 0.09789f
C34 uio_oe[1] VGND 0.09789f
C35 uio_oe[2] VGND 0.09789f
C36 uio_oe[3] VGND 0.09789f
C37 uio_oe[4] VGND 0.09789f
C38 uio_oe[5] VGND 0.09789f
C39 uio_oe[6] VGND 0.09789f
C40 uio_oe[7] VGND 0.09789f
C41 ua[1] VGND 23.692f
C42 ui_in[1] VGND 36.1476f
C43 ui_in[0] VGND 34.1105f
C44 ua[2] VGND 26.9787f
C45 ua[3] VGND 30.6744f
C46 ui_in[3] VGND 22.8547f
C47 ua[0] VGND 87.9149f
C48 ui_in[4] VGND 35.4304f
C49 ui_in[2] VGND 20.4959f
C50 ua[4] VGND 33.8355f
C51 VDPWR VGND 1.2125p
C52 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VGND 11.5065f
C53 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VGND 4.48926f
C54 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VGND 2.83622f
C55 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_136 VGND 1.22562f
C56 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_135 VGND 1.22562f
C57 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_134 VGND 1.22562f
C58 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_133 VGND 1.22629f
C59 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_132 VGND 1.22562f
C60 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_131 VGND 1.22762f
C61 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_130 VGND 1.22562f
C62 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_129 VGND 1.22562f
C63 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_128 VGND 1.22629f
C64 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_127 VGND 1.22696f
C65 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_126 VGND 1.22562f
C66 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_125 VGND 1.22562f
C67 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_124 VGND 1.22562f
C68 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_123 VGND 1.22629f
C69 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_122 VGND 1.22696f
C70 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_121 VGND 1.22762f
C71 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_120 VGND 1.22562f
C72 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_119 VGND 1.22562f
C73 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_118 VGND 1.22562f
C74 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_117 VGND 1.22696f
C75 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_116 VGND 1.22562f
C76 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_115 VGND 1.22562f
C77 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_114 VGND 1.22562f
C78 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_113 VGND 1.22629f
C79 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_112 VGND 1.22562f
C80 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_111 VGND 1.22762f
C81 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_110 VGND 1.22562f
C82 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_109 VGND 1.22562f
C83 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_108 VGND 1.22629f
C84 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_107 VGND 1.22696f
C85 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_106 VGND 1.22762f
C86 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_105 VGND 1.22562f
C87 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_104 VGND 1.22562f
C88 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_103 VGND 1.22629f
C89 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_102 VGND 1.22696f
C90 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_101 VGND 1.22762f
C91 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_100 VGND 1.22562f
C92 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_98 VGND 1.22629f
C93 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_97 VGND 1.22696f
C94 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_96 VGND 1.22562f
C95 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_95 VGND 1.22562f
C96 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_94 VGND 1.22562f
C97 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_93 VGND 1.22629f
C98 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_92 VGND 1.22696f
C99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_91 VGND 1.22762f
C100 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_90 VGND 1.22562f
C101 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_89 VGND 1.22562f
C102 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_88 VGND 1.22562f
C103 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_87 VGND 1.22696f
C104 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_86 VGND 1.22562f
C105 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_85 VGND 1.22562f
C106 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_84 VGND 1.22562f
C107 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_83 VGND 1.22629f
C108 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_82 VGND 1.22696f
C109 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_81 VGND 1.22762f
C110 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_80 VGND 1.22562f
C111 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_79 VGND 1.22562f
C112 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_78 VGND 1.22629f
C113 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_77 VGND 1.22696f
C114 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_76 VGND 1.22562f
C115 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_75 VGND 1.22562f
C116 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_74 VGND 1.22562f
C117 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_73 VGND 1.22629f
C118 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_72 VGND 1.22696f
C119 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_71 VGND 1.22562f
C120 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_70 VGND 1.22562f
C121 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_69 VGND 1.22562f
C122 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_68 VGND 1.22629f
C123 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_67 VGND 1.22696f
C124 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_66 VGND 1.22762f
C125 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_65 VGND 1.22562f
C126 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_64 VGND 1.22562f
C127 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_63 VGND 1.22629f
C128 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_62 VGND 1.22696f
C129 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_61 VGND 1.22762f
C130 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_60 VGND 1.22562f
C131 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_59 VGND 1.22562f
C132 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_58 VGND 1.22629f
C133 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_57 VGND 1.22562f
C134 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_56 VGND 1.22762f
C135 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_55 VGND 1.22562f
C136 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_54 VGND 1.22562f
C137 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_53 VGND 1.22629f
C138 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_52 VGND 1.22696f
C139 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_51 VGND 1.22762f
C140 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_50 VGND 1.22562f
C141 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_49 VGND 1.22562f
C142 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_48 VGND 1.22629f
C143 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_47 VGND 1.22696f
C144 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_46 VGND 1.22562f
C145 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_45 VGND 1.22562f
C146 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_44 VGND 1.22562f
C147 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_43 VGND 1.22629f
C148 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_42 VGND 1.22696f
C149 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_41 VGND 1.22762f
C150 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_40 VGND 1.22562f
C151 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_39 VGND 1.22562f
C152 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_38 VGND 1.22629f
C153 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_37 VGND 1.22696f
C154 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n VGND 56.048f
C155 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_35 VGND 1.22829f
C156 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_34 VGND 1.22562f
C157 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_33 VGND 1.22629f
C158 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_32 VGND 1.22696f
C159 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_31 VGND 1.22762f
C160 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_30 VGND 1.22562f
C161 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_29 VGND 1.22562f
C162 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_28 VGND 1.22629f
C163 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_27 VGND 1.22696f
C164 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_26 VGND 1.22562f
C165 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_25 VGND 1.22562f
C166 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_24 VGND 1.22562f
C167 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_23 VGND 1.22629f
C168 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_22 VGND 1.22696f
C169 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_21 VGND 1.22762f
C170 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_20 VGND 1.22562f
C171 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_19 VGND 1.22562f
C172 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_18 VGND 1.22629f
C173 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n VGND 78.81621f
C174 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_16 VGND 1.22562f
C175 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_15 VGND 1.22562f
C176 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_14 VGND 1.22562f
C177 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_13 VGND 1.22629f
C178 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_12 VGND 1.22562f
C179 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_11 VGND 1.22762f
C180 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_10 VGND 1.22562f
C181 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_9 VGND 1.22562f
C182 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_8 VGND 1.22629f
C183 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_7 VGND 1.22696f
C184 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_6 VGND 1.22562f
C185 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_5 VGND 1.22562f
C186 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_4 VGND 1.22562f
C187 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_3 VGND 1.22629f
C188 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_2 VGND 1.22896f
C189 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_1 VGND 1.22562f
C190 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_0 VGND 1.22562f
C191 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VGND 14.3155f
C192 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VGND 4.48926f
C193 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VGND 7.66312f
C194 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VGND 7.89561f
C195 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin VGND 2.82434f
C196 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C197 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C198 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VGND 2.49069f
C199 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C200 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C201 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C202 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C203 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C204 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VGND 2.49069f
C205 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C206 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C207 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VGND 11.5086f
C208 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VGND 4.48926f
C209 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VGND 2.83622f
C210 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C211 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C212 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VGND 5.82216f
C213 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C214 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND 51.5669f
C215 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C216 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C217 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND 71.3916f
C218 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C219 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C220 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VGND 5.82216f
C221 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C222 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 VGND 33.3927f
C223 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND 75.0436f
C224 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C225 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VGND 37.237f
C226 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VGND 14.3155f
C227 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VGND 4.48926f
C228 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VGND 7.66312f
C229 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VGND 7.89561f
C230 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin VGND 2.82434f
C231 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND 77.9315f
C232 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_136 VGND 1.22562f
C233 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_135 VGND 1.22562f
C234 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_134 VGND 1.22562f
C235 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_133 VGND 1.22562f
C236 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_132 VGND 1.22696f
C237 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_131 VGND 1.22562f
C238 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_130 VGND 1.22562f
C239 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_129 VGND 1.22562f
C240 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_128 VGND 1.22629f
C241 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_127 VGND 1.22562f
C242 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_126 VGND 1.22562f
C243 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_125 VGND 1.22562f
C244 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_124 VGND 1.22562f
C245 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_123 VGND 1.22629f
C246 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_122 VGND 1.22696f
C247 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_121 VGND 1.22562f
C248 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_120 VGND 1.22562f
C249 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_119 VGND 1.22629f
C250 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_118 VGND 1.22629f
C251 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_117 VGND 1.22562f
C252 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_116 VGND 1.22562f
C253 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_115 VGND 1.22562f
C254 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_114 VGND 1.22562f
C255 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_113 VGND 1.22562f
C256 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_112 VGND 1.22696f
C257 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_111 VGND 1.22562f
C258 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_110 VGND 1.22562f
C259 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_109 VGND 1.22562f
C260 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_108 VGND 1.22629f
C261 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_107 VGND 1.22696f
C262 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_106 VGND 1.22562f
C263 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_105 VGND 1.22562f
C264 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_104 VGND 1.22562f
C265 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_103 VGND 1.22629f
C266 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_102 VGND 1.22696f
C267 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_101 VGND 1.22562f
C268 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_100 VGND 1.22562f
C269 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 VGND 39.0581f
C270 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_98 VGND 1.22629f
C271 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_97 VGND 1.22562f
C272 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_96 VGND 1.22562f
C273 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_95 VGND 1.22562f
C274 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_94 VGND 1.22562f
C275 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_93 VGND 1.22629f
C276 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_92 VGND 1.22696f
C277 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_91 VGND 1.22562f
C278 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_90 VGND 1.22562f
C279 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_89 VGND 1.22629f
C280 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_88 VGND 1.22629f
C281 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_87 VGND 1.22562f
C282 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_86 VGND 1.22562f
C283 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_85 VGND 1.22562f
C284 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_84 VGND 1.22562f
C285 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_83 VGND 1.22629f
C286 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_82 VGND 1.22696f
C287 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_81 VGND 1.22562f
C288 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_80 VGND 1.22562f
C289 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_79 VGND 1.22562f
C290 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_78 VGND 1.22629f
C291 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_77 VGND 1.22562f
C292 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_76 VGND 1.22562f
C293 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_75 VGND 1.22562f
C294 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_74 VGND 1.22562f
C295 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_73 VGND 1.22629f
C296 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_72 VGND 1.22562f
C297 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_71 VGND 1.22562f
C298 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_70 VGND 1.22562f
C299 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_69 VGND 1.22562f
C300 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_68 VGND 1.22629f
C301 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_67 VGND 1.22696f
C302 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_66 VGND 1.22562f
C303 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_65 VGND 1.22562f
C304 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_64 VGND 1.22562f
C305 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_63 VGND 1.22629f
C306 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_62 VGND 1.22696f
C307 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_61 VGND 1.22562f
C308 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_60 VGND 1.22562f
C309 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_59 VGND 1.22562f
C310 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_58 VGND 1.22562f
C311 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_57 VGND 1.22696f
C312 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_56 VGND 1.22562f
C313 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_55 VGND 1.22562f
C314 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_54 VGND 1.22562f
C315 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_53 VGND 1.22629f
C316 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_52 VGND 1.22696f
C317 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_51 VGND 1.22562f
C318 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_50 VGND 1.22562f
C319 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_49 VGND 1.22562f
C320 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_48 VGND 1.22629f
C321 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_47 VGND 1.22562f
C322 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_46 VGND 1.22562f
C323 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_45 VGND 1.22562f
C324 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_44 VGND 1.22562f
C325 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_43 VGND 1.22629f
C326 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_42 VGND 1.22696f
C327 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_41 VGND 1.22562f
C328 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_40 VGND 1.22562f
C329 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_39 VGND 1.22562f
C330 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_38 VGND 1.22629f
C331 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_37 VGND 1.22562f
C332 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p VGND 59.6624f
C333 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_35 VGND 1.22562f
C334 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_34 VGND 1.22562f
C335 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_33 VGND 1.22629f
C336 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_32 VGND 1.22696f
C337 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_31 VGND 1.22562f
C338 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_30 VGND 1.22562f
C339 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_29 VGND 1.22562f
C340 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_28 VGND 1.22629f
C341 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_27 VGND 1.22562f
C342 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_26 VGND 1.22562f
C343 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_25 VGND 1.22562f
C344 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_24 VGND 1.22562f
C345 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_23 VGND 1.22629f
C346 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_22 VGND 1.22696f
C347 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_21 VGND 1.22562f
C348 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_20 VGND 1.22562f
C349 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_19 VGND 1.22562f
C350 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_18 VGND 1.22629f
C351 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p VGND 80.2351f
C352 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_16 VGND 1.22562f
C353 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_15 VGND 1.22562f
C354 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_14 VGND 1.22562f
C355 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_13 VGND 1.22562f
C356 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_12 VGND 1.22696f
C357 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_11 VGND 1.22562f
C358 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_10 VGND 1.22562f
C359 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_9 VGND 1.22562f
C360 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_8 VGND 1.22629f
C361 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_7 VGND 1.22562f
C362 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_6 VGND 1.22562f
C363 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_5 VGND 1.22562f
C364 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_4 VGND 1.22562f
C365 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_3 VGND 1.22896f
C366 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_2 VGND 1.22562f
C367 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_1 VGND 1.22562f
C368 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_0 VGND 1.22562f
C369 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VGND 11.5065f
C370 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VGND 4.48926f
C371 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VGND 2.83622f
C372 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_136 VGND 1.22562f
C373 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_135 VGND 1.22562f
C374 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_134 VGND 1.22562f
C375 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_133 VGND 1.22629f
C376 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_132 VGND 1.22562f
C377 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_131 VGND 1.22762f
C378 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_130 VGND 1.22562f
C379 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_129 VGND 1.22562f
C380 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_128 VGND 1.22629f
C381 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_127 VGND 1.22696f
C382 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_126 VGND 1.22562f
C383 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_125 VGND 1.22562f
C384 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_124 VGND 1.22562f
C385 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_123 VGND 1.22629f
C386 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_122 VGND 1.22696f
C387 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_121 VGND 1.22762f
C388 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_120 VGND 1.22562f
C389 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_119 VGND 1.22562f
C390 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_118 VGND 1.22562f
C391 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_117 VGND 1.22696f
C392 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_116 VGND 1.22562f
C393 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_115 VGND 1.22562f
C394 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_114 VGND 1.22562f
C395 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_113 VGND 1.22629f
C396 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_112 VGND 1.22562f
C397 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_111 VGND 1.22762f
C398 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_110 VGND 1.22562f
C399 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_109 VGND 1.22562f
C400 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_108 VGND 1.22629f
C401 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_107 VGND 1.22696f
C402 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_106 VGND 1.22762f
C403 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_105 VGND 1.22562f
C404 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_104 VGND 1.22562f
C405 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_103 VGND 1.22629f
C406 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_102 VGND 1.22696f
C407 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_101 VGND 1.22762f
C408 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_100 VGND 1.22562f
C409 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_98 VGND 1.22629f
C410 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_97 VGND 1.22696f
C411 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_96 VGND 1.22562f
C412 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_95 VGND 1.22562f
C413 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_94 VGND 1.22562f
C414 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_93 VGND 1.22629f
C415 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_92 VGND 1.22696f
C416 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_91 VGND 1.22762f
C417 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_90 VGND 1.22562f
C418 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_89 VGND 1.22562f
C419 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_88 VGND 1.22562f
C420 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_87 VGND 1.22696f
C421 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_86 VGND 1.22562f
C422 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_85 VGND 1.22562f
C423 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_84 VGND 1.22562f
C424 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_83 VGND 1.22629f
C425 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_82 VGND 1.22696f
C426 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_81 VGND 1.22762f
C427 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_80 VGND 1.22562f
C428 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_79 VGND 1.22562f
C429 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_78 VGND 1.22629f
C430 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_77 VGND 1.22696f
C431 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_76 VGND 1.22562f
C432 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_75 VGND 1.22562f
C433 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_74 VGND 1.22562f
C434 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_73 VGND 1.22629f
C435 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_72 VGND 1.22696f
C436 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_71 VGND 1.22562f
C437 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_70 VGND 1.22562f
C438 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_69 VGND 1.22562f
C439 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_68 VGND 1.22629f
C440 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_67 VGND 1.22696f
C441 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_66 VGND 1.22762f
C442 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_65 VGND 1.22562f
C443 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_64 VGND 1.22562f
C444 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_63 VGND 1.22629f
C445 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_62 VGND 1.22696f
C446 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_61 VGND 1.22762f
C447 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_60 VGND 1.22562f
C448 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_59 VGND 1.22562f
C449 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_58 VGND 1.22629f
C450 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_57 VGND 1.22562f
C451 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_56 VGND 1.22762f
C452 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_55 VGND 1.22562f
C453 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_54 VGND 1.22562f
C454 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_53 VGND 1.22629f
C455 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_52 VGND 1.22696f
C456 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_51 VGND 1.22762f
C457 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_50 VGND 1.22562f
C458 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_49 VGND 1.22562f
C459 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_48 VGND 1.22629f
C460 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_47 VGND 1.22696f
C461 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_46 VGND 1.22562f
C462 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_45 VGND 1.22562f
C463 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_44 VGND 1.22562f
C464 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_43 VGND 1.22629f
C465 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_42 VGND 1.22696f
C466 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_41 VGND 1.22762f
C467 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_40 VGND 1.22562f
C468 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_39 VGND 1.22562f
C469 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_38 VGND 1.22629f
C470 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_37 VGND 1.22696f
C471 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n VGND 59.4865f
C472 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_35 VGND 1.22829f
C473 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_34 VGND 1.22562f
C474 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_33 VGND 1.22629f
C475 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_32 VGND 1.22696f
C476 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_31 VGND 1.22762f
C477 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_30 VGND 1.22562f
C478 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_29 VGND 1.22562f
C479 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_28 VGND 1.22629f
C480 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_27 VGND 1.22696f
C481 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_26 VGND 1.22562f
C482 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_25 VGND 1.22562f
C483 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_24 VGND 1.22562f
C484 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_23 VGND 1.22629f
C485 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_22 VGND 1.22696f
C486 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_21 VGND 1.22762f
C487 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_20 VGND 1.22562f
C488 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_19 VGND 1.22562f
C489 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_18 VGND 1.22629f
C490 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n VGND 79.4888f
C491 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_16 VGND 1.22562f
C492 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_15 VGND 1.22562f
C493 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_14 VGND 1.22562f
C494 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_13 VGND 1.22629f
C495 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_12 VGND 1.22562f
C496 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_11 VGND 1.22762f
C497 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_10 VGND 1.22562f
C498 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_9 VGND 1.22562f
C499 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_8 VGND 1.22629f
C500 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_7 VGND 1.22696f
C501 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_6 VGND 1.22562f
C502 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_5 VGND 1.22562f
C503 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_4 VGND 1.22562f
C504 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_3 VGND 1.22629f
C505 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_2 VGND 1.22896f
C506 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_1 VGND 1.22562f
C507 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_0 VGND 1.22562f
C508 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VGND 14.3155f
C509 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VGND 4.48926f
C510 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VGND 7.66312f
C511 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VGND 7.89561f
C512 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin VGND 2.82434f
C513 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C514 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C515 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VGND 2.49069f
C516 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C517 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C518 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C519 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C520 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C521 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VGND 2.49069f
C522 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C523 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C524 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VGND 11.5086f
C525 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VGND 4.48926f
C526 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VGND 2.83622f
C527 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C528 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C529 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VGND 5.82216f
C530 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C531 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND 51.5669f
C532 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C533 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C534 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND 74.2324f
C535 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C536 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C537 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VGND 5.82216f
C538 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C539 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 VGND 36.4777f
C540 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND 75.0436f
C541 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C542 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VGND 37.237f
C543 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VGND 14.3155f
C544 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VGND 4.48926f
C545 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VGND 7.66312f
C546 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VGND 7.89561f
C547 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin VGND 2.82434f
C548 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND 74.9539f
C549 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_136 VGND 1.22562f
C550 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_135 VGND 1.22562f
C551 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_134 VGND 1.22562f
C552 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_133 VGND 1.22562f
C553 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_132 VGND 1.22696f
C554 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_131 VGND 1.22562f
C555 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_130 VGND 1.22562f
C556 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_129 VGND 1.22562f
C557 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_128 VGND 1.22629f
C558 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_127 VGND 1.22562f
C559 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_126 VGND 1.22562f
C560 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_125 VGND 1.22562f
C561 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_124 VGND 1.22562f
C562 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_123 VGND 1.22629f
C563 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_122 VGND 1.22696f
C564 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_121 VGND 1.22562f
C565 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_120 VGND 1.22562f
C566 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_119 VGND 1.22629f
C567 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_118 VGND 1.22629f
C568 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_117 VGND 1.22562f
C569 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_116 VGND 1.22562f
C570 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_115 VGND 1.22562f
C571 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_114 VGND 1.22562f
C572 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_113 VGND 1.22562f
C573 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_112 VGND 1.22696f
C574 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_111 VGND 1.22562f
C575 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_110 VGND 1.22562f
C576 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_109 VGND 1.22562f
C577 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_108 VGND 1.22629f
C578 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_107 VGND 1.22696f
C579 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_106 VGND 1.22562f
C580 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_105 VGND 1.22562f
C581 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_104 VGND 1.22562f
C582 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_103 VGND 1.22629f
C583 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_102 VGND 1.22696f
C584 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_101 VGND 1.22562f
C585 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_100 VGND 1.22562f
C586 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 VGND 36.1864f
C587 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_98 VGND 1.22629f
C588 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_97 VGND 1.22562f
C589 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_96 VGND 1.22562f
C590 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_95 VGND 1.22562f
C591 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_94 VGND 1.22562f
C592 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_93 VGND 1.22629f
C593 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_92 VGND 1.22696f
C594 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_91 VGND 1.22562f
C595 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_90 VGND 1.22562f
C596 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_89 VGND 1.22629f
C597 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_88 VGND 1.22629f
C598 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_87 VGND 1.22562f
C599 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_86 VGND 1.22562f
C600 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_85 VGND 1.22562f
C601 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_84 VGND 1.22562f
C602 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_83 VGND 1.22629f
C603 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_82 VGND 1.22696f
C604 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_81 VGND 1.22562f
C605 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_80 VGND 1.22562f
C606 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_79 VGND 1.22562f
C607 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_78 VGND 1.22629f
C608 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_77 VGND 1.22562f
C609 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_76 VGND 1.22562f
C610 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_75 VGND 1.22562f
C611 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_74 VGND 1.22562f
C612 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_73 VGND 1.22629f
C613 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_72 VGND 1.22562f
C614 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_71 VGND 1.22562f
C615 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_70 VGND 1.22562f
C616 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_69 VGND 1.22562f
C617 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_68 VGND 1.22629f
C618 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_67 VGND 1.22696f
C619 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_66 VGND 1.22562f
C620 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_65 VGND 1.22562f
C621 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_64 VGND 1.22562f
C622 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_63 VGND 1.22629f
C623 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_62 VGND 1.22696f
C624 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_61 VGND 1.22562f
C625 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_60 VGND 1.22562f
C626 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_59 VGND 1.22562f
C627 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_58 VGND 1.22562f
C628 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_57 VGND 1.22696f
C629 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_56 VGND 1.22562f
C630 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_55 VGND 1.22562f
C631 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_54 VGND 1.22562f
C632 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_53 VGND 1.22629f
C633 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_52 VGND 1.22696f
C634 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_51 VGND 1.22562f
C635 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_50 VGND 1.22562f
C636 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_49 VGND 1.22562f
C637 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_48 VGND 1.22629f
C638 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_47 VGND 1.22562f
C639 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_46 VGND 1.22562f
C640 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_45 VGND 1.22562f
C641 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_44 VGND 1.22562f
C642 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_43 VGND 1.22629f
C643 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_42 VGND 1.22696f
C644 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_41 VGND 1.22562f
C645 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_40 VGND 1.22562f
C646 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_39 VGND 1.22562f
C647 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_38 VGND 1.22629f
C648 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_37 VGND 1.22562f
C649 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p VGND 56.026f
C650 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_35 VGND 1.22562f
C651 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_34 VGND 1.22562f
C652 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_33 VGND 1.22629f
C653 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_32 VGND 1.22696f
C654 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_31 VGND 1.22562f
C655 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_30 VGND 1.22562f
C656 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_29 VGND 1.22562f
C657 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_28 VGND 1.22629f
C658 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_27 VGND 1.22562f
C659 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_26 VGND 1.22562f
C660 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_25 VGND 1.22562f
C661 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_24 VGND 1.22562f
C662 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_23 VGND 1.22629f
C663 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_22 VGND 1.22696f
C664 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_21 VGND 1.22562f
C665 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_20 VGND 1.22562f
C666 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_19 VGND 1.22562f
C667 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_18 VGND 1.22629f
C668 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p VGND 78.8372f
C669 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_16 VGND 1.22562f
C670 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_15 VGND 1.22562f
C671 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_14 VGND 1.22562f
C672 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_13 VGND 1.22562f
C673 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_12 VGND 1.22696f
C674 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_11 VGND 1.22562f
C675 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_10 VGND 1.22562f
C676 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_9 VGND 1.22562f
C677 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_8 VGND 1.22629f
C678 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_7 VGND 1.22562f
C679 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_6 VGND 1.22562f
C680 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_5 VGND 1.22562f
C681 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_4 VGND 1.22562f
C682 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_3 VGND 1.22896f
C683 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_2 VGND 1.22562f
C684 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_1 VGND 1.22562f
C685 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_0 VGND 1.22562f
.ends

