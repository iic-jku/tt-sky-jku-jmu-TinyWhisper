magic
tech sky130A
magscale 1 2
timestamp 1761868878
<< metal1 >>
rect -5165 5620 25055 5770
rect -5165 3060 -5115 3170
rect -3075 3155 -2965 3170
rect -3075 3075 -3060 3155
rect -2980 3075 -2965 3155
rect -3075 3060 -2965 3075
rect -410 3155 -300 3170
rect -410 3075 -395 3155
rect -315 3075 -300 3155
rect -410 3060 -300 3075
rect 2255 3155 2365 3170
rect 2255 3075 2270 3155
rect 2350 3075 2365 3155
rect 2255 3060 2365 3075
rect 4405 3155 4515 3170
rect 4405 3075 4420 3155
rect 4500 3075 4515 3155
rect 3040 3065 3780 3070
rect 4405 3060 4515 3075
rect 7070 3155 7180 3170
rect 7070 3075 7085 3155
rect 7165 3075 7180 3155
rect 7070 3060 7180 3075
rect 9735 3155 9845 3170
rect 9735 3075 9750 3155
rect 9835 3075 9845 3155
rect 9735 3060 9845 3075
rect 12400 3155 12510 3170
rect 12400 3075 12415 3155
rect 12495 3075 12510 3155
rect 12400 3060 12510 3075
rect 15065 3155 15175 3170
rect 15065 3075 15080 3155
rect 15160 3075 15175 3155
rect 15065 3060 15175 3075
rect 17730 3155 17840 3170
rect 17730 3075 17745 3155
rect 17825 3075 17840 3155
rect 19880 3155 19990 3170
rect 17730 3060 17840 3075
rect 19880 3075 19895 3155
rect 19975 3075 19990 3155
rect 19880 3060 19990 3075
rect 22545 3155 22655 3170
rect 22545 3075 22560 3155
rect 22640 3075 22655 3155
rect 22545 3060 22655 3075
rect -5165 1680 25055 1830
<< via1 >>
rect -3060 3075 -2980 3155
rect -395 3075 -315 3155
rect 2270 3075 2350 3155
rect 3035 3070 3785 3160
rect 4420 3075 4500 3155
rect 7085 3075 7165 3155
rect 9750 3075 9835 3155
rect 12415 3075 12495 3155
rect 15080 3075 15160 3155
rect 17745 3075 17825 3155
rect 18515 3065 19255 3130
rect 19895 3075 19975 3155
rect 22560 3075 22640 3155
<< metal2 >>
rect -3195 5375 24850 5525
rect -3195 3170 -3110 5375
rect -530 4330 -445 4340
rect -530 4265 -520 4330
rect -455 4265 -445 4330
rect -3225 3060 -3110 3170
rect -3075 3155 -2965 3170
rect -3075 3075 -3060 3155
rect -2980 3075 -2965 3155
rect -3075 3060 -2965 3075
rect -530 3060 -445 4265
rect 2135 4330 2220 4340
rect 2135 4265 2145 4330
rect 2210 4265 2220 4330
rect 2135 3170 2220 4265
rect 6950 4330 7035 4340
rect 6950 4265 6960 4330
rect 7025 4265 7035 4330
rect 6950 3170 7035 4265
rect 12280 4330 12365 4340
rect 12280 4265 12290 4330
rect 12355 4265 12365 4330
rect -410 3155 -300 3170
rect -410 3075 -395 3155
rect -315 3075 -300 3155
rect -410 3060 -300 3075
rect 2135 3155 2365 3170
rect 2135 3075 2270 3155
rect 2350 3075 2365 3155
rect 2135 3060 2365 3075
rect 4255 3060 4365 3170
rect 4405 3155 4515 3170
rect 4405 3075 4420 3155
rect 4500 3075 4515 3155
rect 4405 3060 4515 3075
rect 6915 3060 7035 3170
rect 7070 3155 7180 3170
rect 7070 3075 7085 3155
rect 7165 3075 7180 3155
rect 7070 3060 7180 3075
rect 4280 2980 4365 3060
rect 4280 2915 4290 2980
rect 4355 2915 4365 2980
rect 4280 2905 4365 2915
rect 9615 2620 9700 3170
rect 9735 3155 9845 3170
rect 9735 3075 9750 3155
rect 9835 3075 9845 3155
rect 9735 3060 9845 3075
rect 12280 3060 12365 4265
rect 22425 4330 22510 4340
rect 22425 4265 22435 4330
rect 22500 4265 22510 4330
rect 17610 3520 17695 3530
rect 17610 3455 17620 3520
rect 17685 3455 17695 3520
rect 12400 3155 12510 3170
rect 12400 3075 12415 3155
rect 12495 3075 12510 3155
rect 12400 3060 12510 3075
rect 9615 2555 9625 2620
rect 9690 2555 9700 2620
rect 9615 2545 9700 2555
rect 14945 2610 15030 3170
rect 15065 3155 15175 3170
rect 15065 3075 15080 3155
rect 15160 3075 15175 3155
rect 15065 3060 15175 3075
rect 17610 3060 17695 3455
rect 22425 3170 22510 4265
rect 25090 4330 25175 4340
rect 25090 4265 25100 4330
rect 25165 4265 25175 4330
rect 17730 3155 17840 3170
rect 17730 3075 17745 3155
rect 17825 3075 17840 3155
rect 19880 3155 19990 3170
rect 17730 3060 17840 3075
rect 19880 3075 19895 3155
rect 19975 3075 19990 3155
rect 19880 3060 19990 3075
rect 22300 3160 22510 3170
rect 22300 3070 22310 3160
rect 22415 3070 22510 3160
rect 22300 3060 22510 3070
rect 22545 3155 22655 3170
rect 22545 3075 22560 3155
rect 22640 3075 22655 3155
rect 22545 3060 22655 3075
rect 25090 3060 25175 4265
rect 14945 2545 14955 2610
rect 15020 2545 15030 2610
rect 14945 2535 15030 2545
<< via2 >>
rect -520 4265 -455 4330
rect -3060 3075 -2980 3155
rect 2145 4265 2210 4330
rect 6960 4265 7025 4330
rect 12290 4265 12355 4330
rect -395 3075 -315 3155
rect 4420 3075 4500 3155
rect 7085 3075 7165 3155
rect 4290 2915 4355 2980
rect 9750 3075 9835 3155
rect 22435 4265 22500 4330
rect 17620 3455 17685 3520
rect 12415 3075 12495 3155
rect 9625 2555 9690 2620
rect 15080 3075 15160 3155
rect 25100 4265 25165 4330
rect 17745 3075 17825 3155
rect 19895 3075 19975 3155
rect 22310 3070 22415 3160
rect 22560 3075 22640 3155
rect 14955 2545 15020 2610
<< metal3 >>
rect -5165 5525 4480 5620
rect -3085 3170 -3000 5525
rect -530 4330 2220 4340
rect -530 4265 -520 4330
rect -455 4265 2145 4330
rect 2210 4265 2220 4330
rect -530 4255 2220 4265
rect 4395 3170 4480 5525
rect 6950 5525 25090 5620
rect 6950 4330 7035 5525
rect 6950 4265 6960 4330
rect 7025 4265 7035 4330
rect 6950 4255 7035 4265
rect 12280 4330 12365 5525
rect 12280 4265 12290 4330
rect 12355 4265 12365 4330
rect 12280 4255 12365 4265
rect 5670 3520 17695 3530
rect 5670 3455 17620 3520
rect 17685 3455 17695 3520
rect 5670 3445 17695 3455
rect -3085 3155 -2965 3170
rect -3085 3075 -3060 3155
rect -2980 3075 -2965 3155
rect -3085 3060 -2965 3075
rect -420 3155 -300 3170
rect -420 3075 -395 3155
rect -315 3075 -300 3155
rect -420 3060 -300 3075
rect 4395 3155 4515 3170
rect 4395 3075 4420 3155
rect 4500 3075 4515 3155
rect 4395 3060 4515 3075
rect -420 1925 -335 3060
rect 4280 2980 4365 2990
rect 4280 2915 4290 2980
rect 4355 2915 4365 2980
rect 4280 2785 4365 2915
rect 5670 2785 5760 3445
rect 9725 3170 9810 3445
rect 12390 3170 12475 3445
rect 19870 3170 19955 5525
rect 22425 4330 25175 4340
rect 22425 4265 22435 4330
rect 22500 4265 25100 4330
rect 25165 4265 25175 4330
rect 22425 4255 25175 4265
rect 4280 2700 5760 2785
rect 7060 3155 7180 3170
rect 7060 3075 7085 3155
rect 7165 3075 7180 3155
rect 7060 3060 7180 3075
rect 9725 3155 9845 3170
rect 9725 3075 9750 3155
rect 9835 3075 9845 3155
rect 9725 3060 9845 3075
rect 12390 3155 12510 3170
rect 12390 3075 12415 3155
rect 12495 3075 12510 3155
rect 12390 3060 12510 3075
rect 15055 3155 15175 3170
rect 15055 3075 15080 3155
rect 15160 3075 15175 3155
rect 15055 3060 15175 3075
rect 17720 3155 17840 3170
rect 17720 3075 17745 3155
rect 17825 3075 17840 3155
rect 17720 3060 17840 3075
rect 19870 3155 19990 3170
rect 19870 3075 19895 3155
rect 19975 3075 19990 3155
rect 19870 3060 19990 3075
rect 21145 3160 22425 3170
rect 21145 3070 22310 3160
rect 22415 3070 22425 3160
rect 21145 3060 22425 3070
rect 22535 3155 22655 3170
rect 22535 3075 22560 3155
rect 22640 3075 22655 3155
rect 22535 3060 22655 3075
rect 7060 1925 7145 3060
rect 15055 2785 15140 3060
rect 17720 2785 17805 3060
rect 21145 2785 21235 3060
rect 15055 2700 21235 2785
rect -5165 1830 7145 1925
rect 9615 2620 9700 2630
rect 9615 2555 9625 2620
rect 9690 2555 9700 2620
rect 9615 1925 9700 2555
rect 14945 2610 15030 2620
rect 14945 2545 14955 2610
rect 15020 2545 15030 2610
rect 14945 1925 15030 2545
rect 22535 1925 22620 3060
rect 9615 1830 25090 1925
use inverter_lv_en_NF4  inverter_lv_en_NF4_0 inverter/inverter_lv_en_NF4
timestamp 1757014995
transform 1 0 2495 0 1 1075
box -165 605 1770 4695
use inverter_lv_en_NF4  inverter_lv_en_NF4_1
timestamp 1757014995
transform 1 0 17970 0 1 1075
box -165 605 1770 4695
use inverter_lv_en_NF6  inverter_lv_en_NF6_0 inverter/inverter_lv_en_NF6
timestamp 1761843949
transform 1 0 -2835 0 1 1075
box -165 605 2305 4695
use inverter_lv_en_NF6  inverter_lv_en_NF6_1
timestamp 1761843949
transform 1 0 -170 0 1 1075
box -165 605 2305 4695
use inverter_lv_en_NF6  inverter_lv_en_NF6_2
timestamp 1761843949
transform 1 0 4645 0 1 1075
box -165 605 2305 4695
use inverter_lv_en_NF6  inverter_lv_en_NF6_3
timestamp 1761843949
transform 1 0 7310 0 1 1075
box -165 605 2305 4695
use inverter_lv_en_NF6  inverter_lv_en_NF6_4
timestamp 1761843949
transform 1 0 9975 0 1 1075
box -165 605 2305 4695
use inverter_lv_en_NF6  inverter_lv_en_NF6_5
timestamp 1761843949
transform 1 0 12640 0 1 1075
box -165 605 2305 4695
use inverter_lv_en_NF6  inverter_lv_en_NF6_6
timestamp 1761843949
transform 1 0 15305 0 1 1075
box -165 605 2305 4695
use inverter_lv_en_NF6  inverter_lv_en_NF6_7
timestamp 1761843949
transform 1 0 20120 0 1 1075
box -165 605 2305 4695
use inverter_lv_en_NF6  inverter_lv_en_NF6_8
timestamp 1761843949
transform 1 0 22785 0 1 1075
box -165 605 2305 4695
use inverter_lv_NF4  inverter_lv_NF4_0 inverter/inverter_lv_NF4
timestamp 1757014995
transform 1 0 -4985 0 1 1075
box -165 605 1770 4695
<< labels >>
flabel metal1 -5145 1750 -5145 1750 0 FreeSans 400 0 0 0 VSS
port 3 nsew
flabel metal1 -5150 5695 -5150 5695 0 FreeSans 400 0 0 0 VDD
port 5 nsew
flabel metal2 -2925 5445 -2925 5445 0 FreeSans 320 0 0 0 ota_core_en_n
flabel metal3 -5150 5570 -5150 5570 0 FreeSans 320 0 0 0 vinp
port 11 nsew
flabel metal3 -5145 1875 -5145 1875 0 FreeSans 320 0 0 0 vinn
port 18 nsew
flabel metal1 -5155 3110 -5155 3110 0 FreeSans 320 0 0 0 di_ota_core_en
port 20 nsew
flabel metal3 25075 5570 25075 5570 0 FreeSans 400 0 0 0 voutn
port 26 nsew
flabel metal3 25075 1880 25075 1880 0 FreeSans 400 0 0 0 voutp
port 28 nsew
<< end >>
