magic
tech sky130A
magscale 1 2
timestamp 1762794087
<< locali >>
rect -3545 1065 27010 3705
rect 27610 2805 35650 3690
rect 27610 1070 35650 1955
<< viali >>
rect -4055 7015 -3910 7235
rect -4055 -3685 -3910 -3465
<< metal1 >>
rect -3820 10060 -3545 10465
rect 3785 10460 4010 10470
rect 3785 10065 3795 10460
rect 4000 10065 4010 10460
rect 3785 10055 4010 10065
rect -5600 9770 -3545 9780
rect -5600 9445 -5590 9770
rect -4410 9445 -3545 9770
rect 27400 9740 27520 9890
rect -5600 9435 -3545 9445
rect -4070 7240 -3545 7250
rect -4070 7010 -4060 7240
rect -3905 7010 -3545 7240
rect -4070 7000 -3545 7010
rect 27400 5570 27520 5720
rect -3820 5015 -3545 5420
rect 3785 5235 4010 5240
rect 3785 5025 3795 5235
rect 4000 5025 4010 5235
rect 3785 5015 4010 5025
rect -3545 2050 27010 3710
rect -3545 1735 -3535 2050
rect -2375 1735 27010 2050
rect -3545 1070 27010 1735
rect -3535 735 -2375 1070
rect -3820 -640 -3595 -235
rect -5600 -930 -3545 -920
rect -5600 -1255 -5590 -930
rect -4410 -1255 -3545 -930
rect 27400 -960 27520 -810
rect -5600 -1265 -3545 -1255
rect -4070 -3460 -3560 -3450
rect -4070 -3690 -4060 -3460
rect -3905 -3690 -3560 -3460
rect -4070 -3700 -3560 -3690
rect 27400 -5130 27520 -4980
rect -3820 -5685 -3545 -5280
rect 3785 -5285 4010 -5275
rect 3785 -5680 3795 -5285
rect 4000 -5680 4010 -5285
rect 3785 -5690 4010 -5680
<< via1 >>
rect 3795 10065 4000 10460
rect -5590 9445 -4410 9770
rect -4060 7235 -3905 7240
rect -4060 7015 -4055 7235
rect -4055 7015 -3910 7235
rect -3910 7015 -3905 7235
rect -4060 7010 -3905 7015
rect 3795 5025 4000 5235
rect -3535 1735 -2375 2050
rect -3535 420 -2375 735
rect 3795 -435 4000 -245
rect -5590 -1255 -4410 -930
rect -4060 -3465 -3905 -3460
rect -4060 -3685 -4055 -3465
rect -4055 -3685 -3910 -3465
rect -3910 -3685 -3905 -3465
rect -4060 -3690 -3905 -3685
rect 3795 -5680 4000 -5285
<< metal2 >>
rect 3785 20010 4010 20020
rect 3785 19925 3795 20010
rect 4000 19925 4010 20010
rect 3785 10460 4010 19925
rect 17425 20010 17650 20020
rect 17425 19925 17435 20010
rect 17640 19925 17650 20010
rect 17425 10850 17650 19925
rect 3785 10065 3795 10460
rect 4000 10065 4010 10460
rect 3785 10055 4010 10065
rect -5600 9770 -3590 9780
rect -5600 9445 -5590 9770
rect -4410 9445 -3590 9770
rect -5600 9435 -3590 9445
rect -4070 7240 -3895 7250
rect -4070 7010 -4060 7240
rect -3905 7010 -3895 7240
rect -4070 7000 -3895 7010
rect 3785 5235 4010 5240
rect 3785 5025 3795 5235
rect 4000 5025 4010 5235
rect 3785 5015 4010 5025
rect 17530 4620 22960 4630
rect 17530 4215 22700 4620
rect 22950 4215 22960 4620
rect 17530 4205 22960 4215
rect -3545 2050 -2365 2060
rect -3545 1735 -3535 2050
rect -2375 1735 -2365 2050
rect -3545 735 -2365 1735
rect -3545 420 -3535 735
rect -2375 420 -2365 735
rect -3545 410 -2365 420
rect 17645 555 22960 565
rect 17645 160 22700 555
rect 22950 160 22960 555
rect 17645 150 22960 160
rect 3785 -245 4010 -235
rect 3785 -435 3795 -245
rect 4000 -435 4010 -245
rect 3785 -445 4010 -435
rect -5600 -930 -3590 -920
rect -5600 -1255 -5590 -930
rect -4410 -1255 -3590 -930
rect -5600 -1265 -3590 -1255
rect -4070 -3460 -3895 -3450
rect -4070 -3690 -4060 -3460
rect -3905 -3690 -3895 -3460
rect -4070 -3700 -3895 -3690
rect 3785 -5285 4010 -5275
rect 3785 -5680 3795 -5285
rect 4000 -5680 4010 -5285
rect 3785 -15105 4010 -5680
rect 3785 -15190 3795 -15105
rect 4000 -15190 4010 -15105
rect 3785 -15200 4010 -15190
rect 17425 -15105 17650 -6295
rect 17425 -15190 17435 -15105
rect 17640 -15190 17650 -15105
rect 17425 -15200 17650 -15190
<< via2 >>
rect 3795 19925 4000 20010
rect 17435 19925 17640 20010
rect -5590 9445 -4410 9770
rect -4060 7010 -3905 7240
rect 3795 5025 4000 5235
rect 22700 4215 22950 4620
rect -3535 1735 -2375 2050
rect 22700 160 22950 555
rect 3795 -435 4000 -245
rect -5590 -1255 -4410 -930
rect -4060 -3690 -3905 -3460
rect 3795 -15190 4000 -15105
rect 17435 -15190 17640 -15105
<< metal3 >>
rect 3785 20010 4010 20020
rect 3785 19925 3795 20010
rect 4000 19925 4010 20010
rect 3785 19915 4010 19925
rect 17425 20010 17650 20020
rect 17425 19925 17435 20010
rect 17640 19925 17650 20010
rect 17425 19915 17650 19925
rect 22025 14455 22250 14465
rect 22025 14330 22035 14455
rect 22240 14330 22250 14455
rect 22025 10770 22250 14330
rect 22640 12645 24110 12655
rect 22640 12450 22650 12645
rect 22900 12450 24110 12645
rect 22640 12440 24110 12450
rect 17245 10545 22250 10770
rect 17245 10085 17470 10545
rect -5600 9770 -4400 9780
rect -5600 9445 -5590 9770
rect -4410 9445 -4400 9770
rect -5600 5665 -4400 9445
rect -5600 4500 -5590 5665
rect -4410 4500 -4400 5665
rect -5600 -930 -4400 4500
rect -5600 -1255 -5590 -930
rect -4410 -1255 -4400 -930
rect -5600 -1265 -4400 -1255
rect -4070 7240 -3895 7250
rect -4070 7010 -4060 7240
rect -3905 7010 -3895 7240
rect -4070 -3460 -3895 7010
rect -455 6545 -230 6555
rect -455 6410 -445 6545
rect -240 6410 -230 6545
rect -455 5240 -230 6410
rect 17465 5380 23670 5390
rect -455 5235 4010 5240
rect -455 5025 3795 5235
rect 4000 5025 4010 5235
rect 17465 5055 23410 5380
rect 23660 5055 23670 5380
rect 17465 5045 23670 5055
rect -455 5015 4010 5025
rect 22690 4620 22960 4630
rect 22690 4215 22700 4620
rect 22950 4215 22960 4620
rect 22690 4205 22960 4215
rect 24170 4610 24540 4620
rect 24170 4215 24180 4610
rect 24530 4215 24540 4610
rect 24170 4205 24540 4215
rect -3545 2050 -2365 4040
rect -3545 1735 -3535 2050
rect -2375 1735 -2365 2050
rect -3545 740 -2365 1735
rect 34415 800 34680 7600
rect -3535 735 -2375 740
rect 22690 555 22960 565
rect 22690 160 22700 555
rect 22950 160 22960 555
rect 22690 150 22960 160
rect 24195 555 24565 565
rect 24195 160 24205 555
rect 24555 160 24565 555
rect 24195 150 24565 160
rect -2120 -245 4010 -235
rect -2120 -435 3795 -245
rect 4000 -435 4010 -245
rect -2120 -445 4010 -435
rect 17465 -280 23670 -270
rect -2120 -1690 -1895 -445
rect 17465 -605 23410 -280
rect 23660 -605 23670 -280
rect 35520 -480 36430 4785
rect 17465 -615 23670 -605
rect -2120 -1810 -2110 -1690
rect -1905 -1810 -1895 -1690
rect -2120 -1820 -1895 -1810
rect -4070 -3690 -4060 -3460
rect -3905 -3690 -3895 -3460
rect -4070 -3700 -3895 -3690
rect 17245 -5770 17470 -5310
rect 17245 -5995 22250 -5770
rect 22025 -9555 22250 -5995
rect 22645 -7695 24115 -7685
rect 22645 -7890 22655 -7695
rect 22905 -7890 24115 -7695
rect 22645 -7900 24115 -7890
rect 22025 -9680 22035 -9555
rect 22240 -9680 22250 -9555
rect 22025 -9690 22250 -9680
rect 3785 -15105 4010 -15095
rect 3785 -15190 3795 -15105
rect 4000 -15190 4010 -15105
rect 3785 -15200 4010 -15190
rect 17425 -15105 17650 -15095
rect 17425 -15190 17435 -15105
rect 17640 -15190 17650 -15105
rect 17425 -15200 17650 -15190
<< via3 >>
rect 3795 19925 4000 20010
rect 17435 19925 17640 20010
rect 22035 14330 22240 14455
rect 22650 12450 22900 12645
rect -5590 4500 -4410 5665
rect -445 6410 -240 6545
rect 23410 5055 23660 5380
rect 22700 4215 22950 4620
rect 24180 4215 24530 4610
rect -3535 1735 -2375 2050
rect -3535 420 -2375 735
rect 22700 160 22950 555
rect 24205 160 24555 555
rect 23410 -605 23660 -280
rect -2110 -1810 -1905 -1690
rect 22655 -7890 22905 -7695
rect 22035 -9680 22240 -9555
rect 3795 -15190 4000 -15105
rect 17435 -15190 17640 -15105
<< metal4 >>
rect 2180 19915 3410 20020
rect 15585 19915 16805 20020
rect 22085 14465 22190 14815
rect 23400 14735 23790 14810
rect 22025 14455 22250 14465
rect 22025 14330 22035 14455
rect 22240 14330 22250 14455
rect 22025 14320 22250 14330
rect -455 6545 -230 12705
rect 2815 12600 4045 12705
rect 16225 12600 17445 12705
rect 22640 12645 22910 14605
rect 20670 10795 20940 12600
rect 22640 12450 22650 12645
rect 22900 12450 22910 12645
rect 22640 12440 22910 12450
rect 20670 10525 22960 10795
rect -455 6410 -445 6545
rect -240 6410 -230 6545
rect -455 6400 -230 6410
rect -5600 5665 21610 5675
rect -5600 4500 -5590 5665
rect -4410 4500 21610 5665
rect -5600 4490 21610 4500
rect 22690 4620 22960 10525
rect 23400 5380 23670 14735
rect 23400 5055 23410 5380
rect 23660 5055 23670 5380
rect 23400 5045 23670 5055
rect 24225 4620 24495 14605
rect 22690 4215 22700 4620
rect 22950 4215 22960 4620
rect 22690 4205 22960 4215
rect 24170 4610 24540 4620
rect 24170 4215 24180 4610
rect 24530 4215 24540 4610
rect 24170 4205 24540 4215
rect -3545 2050 -2365 2060
rect -3545 1735 -3535 2050
rect -2375 1735 -2365 2050
rect -3545 735 -2365 1735
rect -3545 420 -3535 735
rect -2375 420 -2365 735
rect -3545 280 -2365 420
rect 22690 555 22960 565
rect -3545 -905 22245 280
rect 22690 160 22700 555
rect 22950 160 22960 555
rect -2120 -1690 -1895 -1680
rect -2120 -1810 -2110 -1690
rect -1905 -1810 -1895 -1690
rect -2120 -7885 -1895 -1810
rect 22690 -5745 22960 160
rect 24195 555 24565 565
rect 24195 160 24205 555
rect 24555 160 24565 555
rect 24195 150 24565 160
rect 20030 -6015 22960 -5745
rect 23400 -280 23670 -270
rect 23400 -605 23410 -280
rect 23660 -605 23670 -280
rect 20030 -7780 20300 -6015
rect 22645 -7695 22915 -7685
rect 2175 -7885 3405 -7780
rect 15585 -7885 16805 -7780
rect 22645 -7890 22655 -7695
rect 22905 -7890 22915 -7695
rect 22025 -9555 22250 -9545
rect 22025 -9680 22035 -9555
rect 22240 -9680 22250 -9555
rect 22025 -9690 22250 -9680
rect 22080 -9785 22195 -9690
rect 22645 -10035 22915 -7890
rect 23400 -9655 23670 -605
rect 23400 -9780 23795 -9655
rect 24245 -10010 24515 150
rect 2820 -15105 4050 -15095
rect 2820 -15190 3795 -15105
rect 4000 -15190 4050 -15105
rect 2820 -15200 4050 -15190
rect 16225 -15105 17445 -15095
rect 16225 -15190 17435 -15105
rect 16225 -15200 17445 -15190
use C1_5x7  C1_5x7_0 /foss/designs/TinyWhisper/magic/iq_modulator/third_order_mfb_lp_filter/capacitors
timestamp 1762704370
transform 1 0 1792 0 1 18970
box -6792 -6370 1032 1050
use C1_5x7  C1_5x7_1
timestamp 1762704370
transform -1 0 4432 0 -1 13650
box -6792 -6370 1032 1050
use C1_5x7  C1_5x7_2
timestamp 1762704370
transform 1 0 1792 0 1 -8830
box -6792 -6370 1032 1050
use C1_5x7  C1_5x7_3
timestamp 1762704370
transform -1 0 4432 0 -1 -14150
box -6792 -6370 1032 1050
use C2_3x7  C2_3x7_0 /foss/designs/TinyWhisper/magic/iq_modulator/third_order_mfb_lp_filter/capacitors
timestamp 1762705970
transform 1 0 18595 0 1 18970
box -6795 -6370 -2365 1050
use C2_3x7  C2_3x7_1
timestamp 1762705970
transform -1 0 14435 0 -1 13650
box -6795 -6370 -2365 1050
use C2_3x7  C2_3x7_2
timestamp 1762705970
transform 1 0 18595 0 1 -8830
box -6795 -6370 -2365 1050
use C2_3x7  C2_3x7_3
timestamp 1762705970
transform -1 0 14435 0 -1 -14150
box -6795 -6370 -2365 1050
use C3_1x5  C3_1x5_0 /foss/designs/TinyWhisper/magic/iq_modulator/third_order_mfb_lp_filter/capacitors
timestamp 1762706219
transform 1 0 21800 0 1 18970
box 0 -4370 1035 1050
use C3_1x5  C3_1x5_1
timestamp 1762706219
transform 1 0 21800 0 1 -10830
box 0 -4370 1035 1050
use C3_1x5  C3_1x5_2
timestamp 1762706219
transform 1 0 23400 0 1 18970
box 0 -4370 1035 1050
use C3_1x5  C3_1x5_3
timestamp 1762706219
transform 1 0 23400 0 1 -10830
box 0 -4370 1035 1050
use decoupling_caps_14x4  decoupling_caps_14x4_0
timestamp 1762702453
transform 1 0 21214 0 1 3545
box -22074 -3370 1032 1050
use iq_modulator_half  iq_modulator_half_0
timestamp 1762793988
transform 1 0 29600 0 1 -765
box -33280 3565 6830 13420
use iq_modulator_half  iq_modulator_half_1
timestamp 1762793988
transform 1 0 29600 0 1 -11465
box -33280 3565 6830 13420
<< labels >>
flabel metal3 35980 1935 35980 1935 0 FreeSans 1600 0 0 0 vout_RF
port 1 nsew
flabel metal1 -3720 5220 -3720 5220 0 FreeSans 1600 0 0 0 vinn_I
port 3 nsew
flabel metal1 -3715 10265 -3715 10265 0 FreeSans 1600 0 0 0 vinp_I
port 5 nsew
flabel metal1 -3700 -440 -3700 -440 0 FreeSans 1600 0 0 0 vinp_Q
port 85 nsew
flabel metal1 -3685 -5485 -3685 -5485 0 FreeSans 1600 0 0 0 vinn_Q
port 87 nsew
flabel metal1 -2865 2545 -2865 2545 0 FreeSans 1600 0 0 0 VSS
port 91 nsew
flabel metal1 -3675 9605 -3675 9605 0 FreeSans 1600 0 0 0 VDD
port 93 nsew
flabel metal1 27460 9815 27460 9815 0 FreeSans 800 0 0 0 di_LO_IX
port 96 nsew
flabel metal1 27460 5650 27460 5650 0 FreeSans 800 0 0 0 di_LO_I
port 98 nsew
flabel metal1 27460 -885 27460 -885 0 FreeSans 800 0 0 0 di_LO_QX
port 100 nsew
flabel metal1 27455 -5055 27455 -5055 0 FreeSans 800 0 0 0 di_LO_Q
port 101 nsew
flabel metal1 -3780 -3595 -3780 -3595 0 FreeSans 1600 0 0 0 di_afe_en
port 110 nsew
<< end >>
