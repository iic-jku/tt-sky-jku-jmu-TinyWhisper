* PEX produced on Mon Nov 10 06:19:26 PM CET 2025 using /foss/tools/sak/iic-pex.sh with m=1 and s=1
* NGSPICE file created from tt_um_TinyWhisper.ext - technology: sky130A

.subckt tt_um_TinyWhisper_pex clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5] ua[6]
+ ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0]
+ uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] VDPWR VGND
X0 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_63 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_64 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_118 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_117 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X2 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X3 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_131 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_132 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X4 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_126 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_125 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X5 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X6 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=279.66 ps=1.9598k w=3 l=0.15
X7 VDPWR ui_in[4] iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X8 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X9 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X10 VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X11 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X12 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X13 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_11 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_12 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X14 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X15 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X16 VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X17 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=173.57899 ps=1.6812k w=1 l=0.15
X18 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X19 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X20 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=29.46 ps=204.67999 w=3 l=0.15
X21 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X22 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_57 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_56 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X23 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_22 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_21 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X24 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_11 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_10 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X25 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X26 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X27 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_65 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_64 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X28 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X29 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X30 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X31 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_10 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_9 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X32 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X33 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X34 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X35 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_34 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_35 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X36 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_20 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_21 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X37 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_63 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_64 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X38 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X39 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X40 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_74 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_75 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X41 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_15 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_14 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X42 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_131 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_132 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X43 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_37 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X44 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_22 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_23 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X45 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_8 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_9 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X46 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X47 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_76 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_77 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X48 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X49 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X50 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_62 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_63 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X51 VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X52 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X53 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_102 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_101 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X54 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_88 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_87 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X55 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_81 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_82 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X56 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=1.27 ps=4.54 w=1 l=0.15
X57 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_90 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_89 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X58 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_76 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_75 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X59 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_130 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_129 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X60 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X61 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=9.82 ps=76.68 w=1 l=0.15
X62 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X63 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X64 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=55.2 ps=372.79999 w=3 l=0.15
X65 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X66 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X67 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X68 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X69 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X70 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_15 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_14 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X71 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X72 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X73 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X74 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X75 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X76 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X77 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_81 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_82 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X78 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X79 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X80 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_26 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_27 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X81 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n ui_in[4] VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X82 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X83 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_52 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_51 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X84 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X85 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=9.82 ps=76.68 w=1 l=0.15
X86 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X87 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X88 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X89 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_40 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_39 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X90 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X91 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X92 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X93 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X94 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=18.4 ps=148.8 w=1 l=0.15
X95 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X96 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X97 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X98 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X99 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X100 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X101 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X102 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X103 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X104 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X105 VGND VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X106 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X107 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X108 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X109 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X110 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X111 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X112 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X113 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X114 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X115 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X116 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X117 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X118 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X119 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X120 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X121 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X122 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X123 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X124 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X125 VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X126 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X127 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X128 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X129 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X130 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X131 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X132 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X133 VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X134 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X135 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X136 VGND VDPWR VGND VGND sky130_fd_pr__pfet_01v8 ad=7.25 pd=50.58 as=511.27039 ps=5.45952k w=25 l=25
X137 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=29.46 ps=204.67999 w=3 l=0.15
X138 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X139 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X140 ui_in[0] VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X141 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X142 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X143 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X144 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=9.82 ps=76.68 w=1 l=0.15
X145 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X146 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X147 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X148 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X149 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X150 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X151 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X152 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X153 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X154 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X155 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X156 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X157 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X158 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X159 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X160 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X161 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X162 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X163 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X164 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X165 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X166 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X167 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X168 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_116 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_115 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X169 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_55 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_56 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X170 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X171 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X172 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_109 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_110 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X173 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X174 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X175 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X176 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_104 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_103 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X177 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X178 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X179 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X180 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_123 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_122 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X181 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_109 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_108 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X182 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=1.27 ps=4.54 w=1 l=0.15
X183 VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X184 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X185 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X186 VGND VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X187 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X188 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X189 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X190 VGND VDPWR sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X191 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X192 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X193 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X194 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X195 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X196 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X197 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_55 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_56 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X198 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X199 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_109 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_110 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X200 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_0 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_1 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X201 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X202 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X203 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X204 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_123 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_122 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X205 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_109 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_108 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X206 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X207 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_59 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_60 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X208 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X209 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_74 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_73 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X210 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X211 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_13 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_14 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X212 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_54 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_53 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X213 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X214 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_128 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_127 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X215 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_122 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_121 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X216 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_67 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_68 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X217 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X218 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X219 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X220 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X221 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_118 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_119 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X222 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_59 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_58 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X223 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_113 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_112 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X224 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X225 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X226 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_120 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_121 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X227 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_135 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_134 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X228 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X229 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_128 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_129 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X230 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X231 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X232 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X233 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X234 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X235 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X236 ui_in[2] VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X237 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X238 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X239 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X240 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=9.82 ps=76.68 w=1 l=0.15
X241 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_59 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_60 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X242 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X243 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X244 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_24 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_25 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X245 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_13 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_14 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X246 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X247 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_67 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_68 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X248 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X249 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X250 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X251 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X252 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X253 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_12 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_13 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X254 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X255 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0 ps=0 w=3 l=1
X256 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_59 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_58 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X257 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_38 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_37 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X258 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_24 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_23 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X259 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_113 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_112 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X260 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_92 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_91 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X261 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_31 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_32 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X262 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_78 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_77 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X263 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_18 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X264 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_135 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_134 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X265 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_3 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_4 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X266 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X267 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_26 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_25 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X268 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X269 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_71 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_72 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X270 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_80 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_79 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X271 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_66 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_65 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X272 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_104 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_105 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X273 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_90 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_91 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X274 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_85 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_84 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X275 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_130 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_131 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X276 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X277 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X278 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_71 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_70 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X279 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_92 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_93 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X280 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X281 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_78 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_79 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X282 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_125 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_124 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X283 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_132 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_133 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X284 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X285 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X286 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X287 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X288 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X289 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_123 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_124 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X290 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X291 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X292 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X293 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X294 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X295 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X296 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X297 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X298 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X299 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X300 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X301 VGND VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X302 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X303 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X304 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_31 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_32 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X305 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_18 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X306 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_3 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_4 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X307 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X308 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X309 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_71 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_72 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X310 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X311 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_2 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_1 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X312 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X313 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X314 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_42 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_41 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X315 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X316 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_28 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_27 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X317 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_85 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_84 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X318 VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X319 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_71 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_70 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X320 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_21 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_22 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X321 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_125 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_124 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X322 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X323 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X324 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_30 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_29 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X325 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_16 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_15 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X326 VGND VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X327 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X328 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_54 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_55 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X329 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X330 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X331 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_40 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_41 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X332 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X333 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X334 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_94 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_95 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X335 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_35 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_34 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X336 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_80 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_81 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X337 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X338 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_21 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_20 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X339 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_42 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_43 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X340 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_123 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_124 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X341 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_28 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_29 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X342 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_96 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_97 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X343 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X344 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X345 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_75 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_74 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X346 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_82 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_83 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X347 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_68 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_69 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X348 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X349 VGND VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X350 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X351 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_108 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_107 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X352 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_94 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_93 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X353 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X354 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_101 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_102 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X355 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_87 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_88 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X356 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_96 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_95 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X357 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X358 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_136 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_135 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X359 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X360 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X361 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X362 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_21 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_22 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X363 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X364 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X365 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_35 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_34 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X366 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_21 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_20 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X367 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X368 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_75 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_74 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X369 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X370 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VGND ui_in[1] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.93 ps=6.62 w=3 l=0.15
X371 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X372 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X373 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X374 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X375 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X376 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_44 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_45 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X377 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_101 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_102 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X378 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X379 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_87 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_88 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X380 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X381 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X382 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_66 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_67 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X383 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_46 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_47 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X384 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_32 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_33 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X385 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X386 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X387 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=29.46 ps=204.67999 w=3 l=0.15
X388 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X389 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_58 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_57 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X390 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X391 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_112 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_111 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X392 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_51 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_52 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X393 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_46 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_45 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X394 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_100 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X395 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X396 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X397 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X398 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X399 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X400 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0 ps=0 w=3 l=1
X401 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X402 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X403 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X404 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X405 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X406 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X407 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X408 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VGND ui_in[3] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.93 ps=6.62 w=3 l=0.15
X409 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X410 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X411 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=0 ps=0 w=9 l=1
X412 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X413 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X414 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X415 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X416 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X417 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X418 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X419 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X420 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X421 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X422 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X423 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X424 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X425 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X426 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X427 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=29.46 ps=204.67999 w=3 l=0.15
X428 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_51 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_52 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X429 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X430 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X431 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_16 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X432 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X433 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X434 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X435 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_2 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_3 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X436 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X437 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X438 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_4 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_5 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X439 VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X440 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X441 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X442 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_70 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_69 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X443 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X444 VGND VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X445 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X446 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X447 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X448 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X449 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X450 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X451 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X452 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_136 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X453 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X454 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X455 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X456 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X457 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X458 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X459 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X460 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X461 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X462 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X463 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X464 VGND VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X465 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X466 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X467 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X468 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X469 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X470 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X471 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X472 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X473 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X474 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X475 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X476 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X477 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X478 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X479 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X480 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X481 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X482 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X483 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X484 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X485 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X486 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=0 ps=0 w=9 l=1
X487 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_115 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_116 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X488 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X489 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X490 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X491 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X492 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X493 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X494 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X495 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X496 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X497 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X498 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X499 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X500 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X501 VGND VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X502 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X503 VGND VDPWR VGND VGND sky130_fd_pr__pfet_01v8 ad=7.25 pd=50.58 as=0 ps=0 w=25 l=25
X504 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X505 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X506 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X507 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X508 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X509 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X510 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X511 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X512 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X513 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=0 ps=0 w=9 l=1
X514 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X515 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X516 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X517 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X518 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X519 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_115 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_116 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X520 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X521 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X522 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X523 VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X524 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X525 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X526 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X527 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X528 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X529 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X530 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X531 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X532 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X533 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X534 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_134 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_133 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X535 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X536 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_73 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_74 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X537 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X538 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X539 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X540 VGND VDPWR VGND VGND sky130_fd_pr__pfet_01v8 ad=7.25 pd=50.58 as=0 ps=0 w=25 l=25
X541 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_127 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_128 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X542 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X543 VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X544 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_119 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_118 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X545 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X546 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X547 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X548 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X549 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X550 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X551 VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X552 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X553 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X554 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X555 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X556 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X557 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X558 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X559 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_30 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_31 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X560 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_73 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_74 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X561 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_25 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_24 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X562 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_127 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_128 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X563 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X564 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_18 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_19 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X565 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X566 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X567 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X568 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_44 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_43 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X569 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X570 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X571 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_119 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_118 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X572 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_98 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_97 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X573 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_37 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_38 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X574 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_84 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_83 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X575 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X576 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_23 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_24 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X577 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X578 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_91 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_92 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X579 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_77 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_78 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X580 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_86 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_85 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X581 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X582 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_110 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_111 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X583 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X584 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X585 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_105 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_104 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X586 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_91 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_90 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X587 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X588 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_98 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X589 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_131 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_130 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X590 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X591 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X592 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X593 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X594 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X595 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X596 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X597 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X598 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_25 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_24 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X599 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X600 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=0 ps=0 w=9 l=1
X601 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X602 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X603 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_37 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_38 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X604 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X605 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X606 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_23 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_24 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X607 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_91 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_92 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X608 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_77 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_78 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X609 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X610 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X611 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X612 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X613 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X614 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_62 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_61 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X615 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_48 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_47 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X616 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X617 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_2 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X618 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_34 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_33 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X619 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_105 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_104 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X620 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_91 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_90 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X621 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X622 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_41 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_42 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X623 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_27 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_28 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X624 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_131 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_130 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X625 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_50 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_49 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X626 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_35 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X627 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X628 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X629 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X630 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X631 VGND VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X632 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_60 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_61 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X633 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X634 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_114 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_115 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X635 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_55 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_54 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X636 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_100 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_101 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X637 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X638 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_41 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_40 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X639 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_48 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_49 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X640 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X641 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X642 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_116 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_117 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X643 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_95 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_94 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X644 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X645 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_102 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_103 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X646 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X647 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_81 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_80 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X648 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X649 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X650 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X651 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_88 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_89 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X652 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X653 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X654 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X655 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_114 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_113 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X656 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_107 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_108 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X657 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_93 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_94 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X658 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X659 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VGND ui_in[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.93 ps=6.62 w=3 l=0.15
X660 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X661 VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X662 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X663 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X664 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_2 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X665 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X666 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X667 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_41 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_42 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X668 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_27 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_28 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X669 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X670 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X671 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_6 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_7 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X672 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X673 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_55 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_54 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X674 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X675 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X676 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_41 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_40 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X677 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X678 VGND VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X679 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_20 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_19 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X680 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_6 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_5 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X681 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_95 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_94 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X682 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_0 ua[4] VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X683 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X684 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X685 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_81 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_80 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X686 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X687 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_8 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_7 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X688 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_50 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_51 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X689 VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X690 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X691 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_107 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_108 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X692 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_86 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_87 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X693 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_93 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_94 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X694 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_72 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_73 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X695 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_45 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_44 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X696 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X697 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X698 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_126 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_127 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X699 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_52 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_53 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X700 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_38 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_39 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X701 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_67 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_66 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X702 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_106 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_107 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X703 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X704 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X705 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_118 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_117 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X706 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X707 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_57 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_58 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X708 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X709 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X710 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X711 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_111 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_112 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X712 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_126 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_125 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X713 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_120 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_119 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X714 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_106 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_105 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X715 VGND VDPWR VGND VGND sky130_fd_pr__pfet_01v8 ad=7.25 pd=50.58 as=0 ps=0 w=25 l=25
X716 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X717 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X718 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X719 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X720 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X721 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X722 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X723 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X724 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X725 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X726 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_45 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_44 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X727 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X728 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X729 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_10 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_9 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X730 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_67 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_66 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X731 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X732 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X733 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X734 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_12 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_11 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X735 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X736 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_57 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_58 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X737 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X738 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X739 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_37 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X740 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_22 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_23 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X741 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_8 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_9 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X742 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_111 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_112 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X743 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X744 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X745 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_76 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_77 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X746 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X747 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_16 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X748 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_62 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_63 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X749 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_56 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_57 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X750 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_3 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_2 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X751 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X752 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_10 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_11 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X753 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X754 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X755 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_64 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_65 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X756 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X757 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X758 VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X759 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X760 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_90 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_89 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X761 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X762 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X763 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_76 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_75 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X764 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X765 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_130 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_129 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X766 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_69 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_70 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X767 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_64 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_63 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X768 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X769 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X770 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_132 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_131 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X771 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X772 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X773 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X774 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X775 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X776 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X777 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X778 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_136 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X779 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X780 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X781 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X782 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X783 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X784 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X785 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X786 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X787 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X788 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X789 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_16 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X790 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_3 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_2 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X791 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X792 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X793 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X794 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_26 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_27 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X795 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X796 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VGND ui_in[2] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.93 ps=6.62 w=3 l=0.15
X797 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X798 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_69 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_70 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X799 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X800 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_14 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_15 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X801 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X802 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X803 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X804 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_40 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_39 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X805 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X806 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin ui_in[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X807 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_136 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X808 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X809 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X810 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_82 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_81 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X811 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X812 VGND VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X813 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X814 VGND VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X815 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X816 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X817 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X818 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n ui_in[4] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X819 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X820 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X821 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X822 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X823 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X824 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=3.81 ps=8.54 w=3 l=0.15
X825 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X826 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X827 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X828 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X829 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X830 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X831 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X832 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X833 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X834 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X835 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X836 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X837 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X838 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X839 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X840 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X841 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X842 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X843 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X844 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X845 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X846 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=3.81 ps=8.54 w=3 l=0.15
X847 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X848 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X849 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X850 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X851 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X852 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X853 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X854 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X855 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X856 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_133 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_134 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X857 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X858 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X859 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X860 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X861 VGND VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X862 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X863 VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X864 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X865 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X866 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=1.27 ps=4.54 w=1 l=0.15
X867 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X868 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X869 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X870 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X871 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X872 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X873 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X874 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X875 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X876 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X877 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X878 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X879 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X880 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X881 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X882 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X883 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X884 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_31 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_30 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X885 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_133 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_134 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X886 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X887 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X888 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X889 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X890 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X891 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X892 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_104 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_103 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X893 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_43 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_44 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X894 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X895 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X896 VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X897 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_97 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_98 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X898 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X899 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_83 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_84 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X900 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X901 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X902 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X903 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X904 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X905 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_111 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_110 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X906 VGND VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X907 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X908 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X909 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_31 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_30 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X910 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X911 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n ui_in[4] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X912 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X913 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X914 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X915 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_0 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_1 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X916 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X917 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X918 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_43 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_44 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X919 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X920 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_97 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_98 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X921 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_83 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_84 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X922 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X923 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X924 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X925 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X926 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X927 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X928 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_54 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_53 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X929 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_111 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_110 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X930 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X931 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_122 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_121 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X932 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_61 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_62 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X933 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_47 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_48 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X934 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X935 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_33 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_34 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X936 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_56 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_55 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X937 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X938 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_110 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_109 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X939 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X940 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X941 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X942 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X943 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X944 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X945 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X946 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_120 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_121 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X947 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_61 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_60 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X948 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X949 VGND VDPWR sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X950 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X951 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_115 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_114 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X952 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_128 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_129 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X953 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X954 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_122 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_123 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X955 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_101 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_100 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X956 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_108 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_109 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X957 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X958 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X959 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X960 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X961 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X962 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X963 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_113 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_114 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X964 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X965 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X966 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X967 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X968 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X969 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X970 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X971 VGND ui_in[2] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X972 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_61 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_62 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X973 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_47 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_48 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X974 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_33 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_34 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X975 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X976 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_12 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_13 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X977 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X978 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_7 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_6 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X979 VGND VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X980 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X981 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X982 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_61 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_60 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X983 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=1.27 ps=4.54 w=1 l=0.15
X984 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_26 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_25 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X985 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_115 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_114 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X986 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_101 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_100 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X987 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_80 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_79 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X988 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_19 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_20 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X989 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_66 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_65 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X990 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_60 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_59 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X991 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_5 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_6 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X992 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X993 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_14 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_13 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X994 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X995 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VDPWR ui_in[1] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X996 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_68 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_67 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X997 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X998 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_113 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_114 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X999 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_92 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_93 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1000 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1001 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_78 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_79 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1002 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_51 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_50 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1003 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_58 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_59 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1004 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_87 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_86 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1005 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1006 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1007 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_132 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_133 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1008 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_73 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_72 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1009 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1010 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_112 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_113 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1011 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_127 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_126 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1012 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1013 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1014 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_134 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_135 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1015 ui_in[1] VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0.495 ps=3.33 w=3 l=0.15
X1016 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1017 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1018 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1019 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1020 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_117 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_118 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1021 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1022 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1023 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1024 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1025 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_125 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_126 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1026 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1027 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_7 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_6 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1028 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1029 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1030 VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X1031 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1032 VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X1033 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_19 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_20 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1034 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_5 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_6 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1035 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1036 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n ui_in[4] VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1037 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1038 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1039 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1040 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_51 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_50 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1041 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_30 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_29 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1042 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_16 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_15 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1043 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_87 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_86 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1044 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1045 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X1046 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_73 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_72 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1047 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1048 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1049 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1050 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_9 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_10 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1051 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_127 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_126 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1052 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_32 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_31 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1053 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1054 ui_in[3] VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0.495 ps=3.33 w=3 l=0.15
X1055 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_18 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1056 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1057 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_4 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_3 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1058 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_72 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_71 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1059 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1060 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1061 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_42 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_43 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1062 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1063 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_28 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_29 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1064 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_117 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_118 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1065 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1066 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin ui_in[0] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1067 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_96 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_97 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1068 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_37 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1069 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1070 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_82 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_83 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1071 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_23 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_22 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1072 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_68 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_69 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1073 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_125 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_126 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1074 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_9 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_8 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1075 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1076 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1077 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_77 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_76 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1078 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_63 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_62 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1079 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_84 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_85 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1080 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_70 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_71 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1081 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_124 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_125 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1082 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1083 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_96 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_95 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1084 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1085 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_89 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_90 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1086 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_136 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_135 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1087 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_75 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_76 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1088 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1089 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1090 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_129 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_130 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1091 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1092 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_124 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_123 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1093 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1094 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1095 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_9 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_10 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1096 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1097 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1098 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1099 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1100 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1101 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1102 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1103 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1104 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin ui_in[2] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1105 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1106 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_37 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1107 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1108 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_23 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_22 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1109 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1110 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_9 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_8 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1111 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_77 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_76 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1112 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1113 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1114 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_63 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_62 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1115 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1116 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_22 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_21 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1117 VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X1118 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1119 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1120 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_46 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_47 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1121 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_32 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_33 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1122 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1123 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_89 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_90 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1124 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_75 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_76 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1125 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1126 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_27 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_26 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1127 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_129 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_130 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1128 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_34 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_35 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1129 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1130 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_20 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_21 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1131 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1132 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1133 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_74 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_75 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1134 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1135 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1136 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_46 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_45 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1137 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_100 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1138 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_39 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_40 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1139 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=3.81 ps=8.54 w=3 l=0.15
X1140 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1141 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1142 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_102 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_101 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1143 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_88 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_87 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1144 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1145 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1146 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1147 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1148 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1149 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1150 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1151 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VDPWR ui_in[3] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X1152 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1153 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1154 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1155 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1156 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1157 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_27 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_26 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1158 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1159 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1160 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1161 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1162 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1163 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1164 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1165 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_39 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_40 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1166 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1167 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1168 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_4 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_5 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1169 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1170 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1171 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1172 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1173 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1174 VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X1175 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1176 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1177 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_52 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_51 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1178 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1179 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n ui_in[4] VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1180 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1181 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=1.27 ps=4.54 w=1 l=0.15
X1182 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1183 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1184 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1185 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1186 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X1187 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1188 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin ui_in[1] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1189 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1190 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1191 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1192 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1193 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1194 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1195 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1196 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1197 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1198 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1199 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X1200 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1201 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1202 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1203 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1204 VGND ui_in[4] iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1205 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1206 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1207 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1208 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1209 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1210 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1211 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1212 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1213 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin ui_in[3] VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1214 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1215 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1216 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1217 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1218 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1219 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1220 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1221 VGND VDPWR VGND VGND sky130_fd_pr__pfet_01v8 ad=7.25 pd=50.58 as=0 ps=0 w=25 l=25
X1222 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1223 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1224 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1225 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1226 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1227 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1228 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1229 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1230 VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X1231 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1232 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin ui_in[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1233 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1234 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1235 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_103 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_104 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1236 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1237 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1238 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1239 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1240 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=3.81 ps=8.54 w=3 l=0.15
X1241 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1242 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1243 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1244 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1245 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1246 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1247 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1248 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1249 VDPWR ui_in[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1250 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1251 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1252 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1253 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1254 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1255 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1256 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1257 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1258 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1259 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_0 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1260 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_103 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_104 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1261 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1262 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_53 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_54 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1263 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_121 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_122 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1264 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1265 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1266 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1267 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_116 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_115 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1268 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1269 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1270 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1271 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1272 VDPWR ui_in[2] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1273 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_121 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_120 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1274 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1275 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_129 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_128 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1276 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1277 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1278 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1279 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=1.27 ps=4.54 w=1 l=0.15
X1280 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1281 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1282 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=1.27 ps=4.54 w=1 l=0.15
X1283 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1284 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_0 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1285 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1286 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1287 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1288 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1289 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1290 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VDPWR ui_in[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X1291 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1292 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1293 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1294 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1295 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1296 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1297 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_53 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_54 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1298 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_121 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_122 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1299 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1300 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_18 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_19 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1301 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X1302 ui_in[0] VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0.495 ps=3.33 w=3 l=0.15
X1303 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1304 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_13 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_12 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1305 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1306 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1307 VGND ui_in[4] iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1308 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1309 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_121 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_120 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1310 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1311 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_86 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_85 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1312 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_25 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_26 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1313 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_129 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_128 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1314 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_79 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_80 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1315 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_65 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_66 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1316 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1317 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_74 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_73 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1318 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1319 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1320 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_128 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_127 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1321 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1322 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1323 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_98 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1324 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1325 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1326 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1327 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1328 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_93 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_92 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1329 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1330 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_79 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_78 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1331 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_118 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_119 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1332 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_133 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_132 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1333 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1334 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1335 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1336 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1337 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1338 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1339 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1340 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1341 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_13 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_12 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1342 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1343 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1344 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1345 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1346 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin ui_in[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1347 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_25 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_26 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1348 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1349 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_79 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_80 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1350 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_65 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_66 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1351 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1352 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1353 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_24 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_25 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1354 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_50 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_49 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1355 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_35 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1356 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_93 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_92 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1357 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_79 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_78 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1358 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1359 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_29 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_30 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1360 VDPWR ui_in[1] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1361 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_133 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_132 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1362 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_38 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_37 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1363 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_15 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_16 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1364 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_24 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_23 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1365 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1366 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_92 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_91 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1367 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_78 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_77 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1368 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1369 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_48 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_49 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1370 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_116 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_117 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1371 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1372 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_102 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_103 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1373 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1374 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1375 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_43 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_42 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1376 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_88 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_89 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1377 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_29 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_28 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1378 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_97 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_96 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1379 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_83 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_82 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1380 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1381 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_104 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_105 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1382 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_69 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_68 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1383 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_90 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_91 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1384 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_130 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_131 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1385 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1386 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1387 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_95 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_96 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1388 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1389 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1390 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_135 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_136 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1391 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X1392 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1393 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1394 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1395 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1396 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1397 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1398 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_29 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_30 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1399 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1400 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_15 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_16 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1401 VDPWR ui_in[3] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1402 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1403 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_0 ua[2] VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1404 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_43 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_42 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1405 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_29 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_28 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1406 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_8 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_7 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1407 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_97 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_96 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1408 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_83 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_82 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1409 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1410 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_2 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_1 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1411 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_69 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_68 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1412 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_42 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_41 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1413 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1414 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_28 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_27 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1415 VGND ui_in[1] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1416 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_52 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_53 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1417 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_38 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_39 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1418 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1419 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_106 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_107 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1420 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_95 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_96 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1421 VDPWR ui_in[4] iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1422 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1423 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_47 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_46 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1424 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1425 VGND VDPWR VGND VGND sky130_fd_pr__pfet_01v8 ad=7.25 pd=50.58 as=0 ps=0 w=25 l=25
X1426 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_54 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_55 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1427 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_33 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_32 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1428 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_135 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_136 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1429 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_40 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_41 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1430 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1431 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VDPWR ui_in[2] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X1432 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1433 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_94 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_95 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1434 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_80 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_81 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1435 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1436 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_120 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_119 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1437 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_106 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_105 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1438 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_45 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_46 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1439 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1440 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_100 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1441 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1442 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1443 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1444 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_108 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_107 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1445 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1446 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_94 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_93 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1447 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1448 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1449 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1450 ui_in[2] VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0.495 ps=3.33 w=3 l=0.15
X1451 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1452 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1453 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1454 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1455 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1456 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1457 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1458 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1459 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1460 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1461 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1462 VGND ui_in[4] iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1463 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1464 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_47 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_46 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1465 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1466 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_33 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_32 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1467 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1468 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_12 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_11 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1469 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1470 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1471 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_45 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_46 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1472 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_56 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_57 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1473 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1474 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_10 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_11 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1475 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_100 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1476 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1477 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_64 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_65 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1478 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1479 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1480 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_5 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_4 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1481 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_44 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_45 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1482 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1483 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1484 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1485 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_66 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_67 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1486 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1487 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1488 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1489 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_64 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_63 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1490 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_58 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_57 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1491 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_132 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_131 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1492 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1493 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_112 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_111 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1494 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1495 VGND VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X1496 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1497 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1498 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1499 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1500 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1501 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_5 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_4 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1502 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1503 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1504 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1505 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1506 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1507 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1508 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1509 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1510 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1511 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1512 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_14 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_15 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1513 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X1514 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_16 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1515 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_2 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_3 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1516 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1517 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin ui_in[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1518 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1519 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1520 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1521 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1522 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1523 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_82 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_81 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1524 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1525 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1526 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1527 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n ui_in[4] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1528 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X1529 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_70 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_69 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1530 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1531 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1532 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1533 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1534 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_136 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1535 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1536 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1537 VGND ui_in[3] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1538 VDPWR ui_in[4] iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1539 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1540 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1541 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1542 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1543 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1544 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=3.81 ps=8.54 w=3 l=0.15
X1545 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1546 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1547 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1548 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1549 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1550 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1551 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1552 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1553 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1554 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1555 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1556 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1557 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1558 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1559 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1560 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1561 VGND VDPWR VGND VGND sky130_fd_pr__pfet_01v8 ad=7.25 pd=50.58 as=0 ps=0 w=25 l=25
X1562 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1563 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1564 VGND ui_in[4] iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1565 VGND VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X1566 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1567 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1568 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1569 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1570 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1571 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=3.81 ps=8.54 w=3 l=0.15
X1572 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1573 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1574 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1575 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1576 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1577 VGND VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X1578 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1579 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1580 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1581 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1582 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1583 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1584 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1585 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1586 VGND VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X1587 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1588 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1589 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1590 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1591 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1592 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1593 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1594 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1595 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1596 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1597 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1598 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_19 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_18 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1599 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1600 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1601 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1602 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_85 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_86 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1603 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_134 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_133 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1604 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1605 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1606 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1607 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_98 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1608 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1609 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1610 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1611 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X1612 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1613 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1614 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n ui_in[4] VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1615 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X1616 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1617 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1618 ui_in[1] VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X1619 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1620 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1621 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1622 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1623 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1624 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1625 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_19 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_18 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1626 VDPWR iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=3.81 ps=8.54 w=3 l=0.15
X1627 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1628 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1629 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1630 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_85 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_86 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1631 VGND VDPWR VGND VGND sky130_fd_pr__pfet_01v8 ad=7.25 pd=50.58 as=0 ps=0 w=25 l=25
X1632 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_30 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_31 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1633 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1634 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1635 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1636 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1637 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_56 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_55 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1638 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1639 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1640 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1641 VDPWR ui_in[4] iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1642 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_110 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_109 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1643 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_98 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1644 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_49 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_50 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1645 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_35 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1646 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1647 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_44 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_43 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1648 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1649 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_98 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_97 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1650 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_84 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_83 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1651 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1652 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_122 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_123 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1653 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1654 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_108 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_109 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1655 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_49 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_48 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1656 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_117 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_116 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1657 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_103 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_102 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1658 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1659 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_89 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_88 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1660 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_110 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_111 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1661 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1662 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1663 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1664 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1665 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1666 VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=3.81 ps=8.54 w=3 l=0.15
X1667 VGND VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X1668 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1669 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1670 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1671 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1672 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1673 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1674 VGND VDPWR iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X1675 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1676 VGND ui_in[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1677 VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X1678 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1679 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_49 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_50 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1680 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_35 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1681 VGND iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=1.27 ps=4.54 w=1 l=0.15
X1682 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n ua[0] VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1683 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1684 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1685 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1686 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1687 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_49 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_48 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1688 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_60 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_59 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1689 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_117 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_116 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1690 ua[1] iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_0 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1691 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_14 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_13 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1692 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_103 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_102 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1693 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_89 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_88 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1694 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_68 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_67 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1695 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_62 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_61 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1696 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_7 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_8 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1697 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_48 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_47 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1698 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_34 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_33 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1699 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1700 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1701 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_58 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_59 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1702 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_112 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_113 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1703 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1704 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1705 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_53 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_52 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1706 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_60 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_61 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1707 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_39 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_38 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1708 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_134 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_135 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1709 ua[0] iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1710 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1711 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_107 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_106 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1712 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1713 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_114 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_115 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1714 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_100 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_101 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1715 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1716 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1717 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_119 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_120 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1718 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_105 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_106 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1719 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1720 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_114 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_113 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1721 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1722 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n ui_in[4] VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1723 VGND iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1724 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1725 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1726 ua[3] iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_0 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1727 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1728 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1729 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1730 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_7 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_8 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1731 VDPWR VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1732 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_6 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_7 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1733 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1734 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl ua[0] VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1735 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_53 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_52 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1736 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_32 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_31 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1737 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_39 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_38 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1738 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDPWR VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1739 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X1740 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_18 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1741 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_107 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_106 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1742 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_4 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_3 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1743 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VDPWR VDPWR sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1744 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_72 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_71 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1745 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_11 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_12 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1746 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_20 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_19 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1747 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1748 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_6 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_5 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1749 ui_in[3] VDPWR iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VGND sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X1750 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1751 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_119 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_120 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1752 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1753 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1754 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_105 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_106 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1755 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1756 VGND VDPWR iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X1757 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_84 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_85 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1758 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_57 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_56 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1759 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_70 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_71 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1760 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_11 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_10 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1761 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_50 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_51 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1762 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1763 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_124 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_125 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1764 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_65 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_64 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1765 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_86 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_87 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1766 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_72 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_73 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1767 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_126 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_127 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1768 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDPWR sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1769 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1770 ua[0] iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1771 VDPWR VGND sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1772 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_124 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_123 VGND sky130_fd_pr__res_xhigh_po_0p35 l=2
X1773 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
C0 ua[5] VGND 0.14696f
C1 ua[6] VGND 0.14696f
C2 ua[7] VGND 0.14696f
C3 ena VGND 0.09789f
C4 clk VGND 0.09789f
C5 rst_n VGND 0.09789f
C6 ui_in[5] VGND 0.09789f
C7 ui_in[6] VGND 0.09789f
C8 ui_in[7] VGND 0.09789f
C9 uio_in[0] VGND 0.09789f
C10 uio_in[1] VGND 0.09789f
C11 uio_in[2] VGND 0.09789f
C12 uio_in[3] VGND 0.09789f
C13 uio_in[4] VGND 0.09789f
C14 uio_in[5] VGND 0.09789f
C15 uio_in[6] VGND 0.09789f
C16 uio_in[7] VGND 0.09789f
C17 ua[1] VGND 23.692f
C18 ui_in[1] VGND 36.1476f
C19 ui_in[0] VGND 34.1105f
C20 ua[2] VGND 26.9787f
C21 ua[3] VGND 30.6744f
C22 ui_in[3] VGND 22.8547f
C23 ua[0] VGND 87.9149f
C24 ui_in[4] VGND 35.4304f
C25 ui_in[2] VGND 20.4959f
C26 ua[4] VGND 33.8355f
C27 VDPWR VGND 1.48787p
C28 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VGND 11.5065f
C29 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VGND 4.48926f
C30 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VGND 2.83622f
C31 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_136 VGND 1.22562f
C32 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_135 VGND 1.22562f
C33 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_134 VGND 1.22562f
C34 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_133 VGND 1.22629f
C35 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_132 VGND 1.22562f
C36 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_131 VGND 1.22762f
C37 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_130 VGND 1.22562f
C38 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_129 VGND 1.22562f
C39 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_128 VGND 1.22629f
C40 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_127 VGND 1.22696f
C41 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_126 VGND 1.22562f
C42 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_125 VGND 1.22562f
C43 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_124 VGND 1.22562f
C44 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_123 VGND 1.22629f
C45 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_122 VGND 1.22696f
C46 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_121 VGND 1.22762f
C47 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_120 VGND 1.22562f
C48 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_119 VGND 1.22562f
C49 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_118 VGND 1.22562f
C50 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_117 VGND 1.22696f
C51 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_116 VGND 1.22562f
C52 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_115 VGND 1.22562f
C53 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_114 VGND 1.22562f
C54 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_113 VGND 1.22629f
C55 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_112 VGND 1.22562f
C56 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_111 VGND 1.22762f
C57 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_110 VGND 1.22562f
C58 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_109 VGND 1.22562f
C59 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_108 VGND 1.22629f
C60 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_107 VGND 1.22696f
C61 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_106 VGND 1.22762f
C62 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_105 VGND 1.22562f
C63 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_104 VGND 1.22562f
C64 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_103 VGND 1.22629f
C65 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_102 VGND 1.22696f
C66 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_101 VGND 1.22762f
C67 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_100 VGND 1.22562f
C68 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_98 VGND 1.22629f
C69 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_97 VGND 1.22696f
C70 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_96 VGND 1.22562f
C71 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_95 VGND 1.22562f
C72 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_94 VGND 1.22562f
C73 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_93 VGND 1.22629f
C74 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_92 VGND 1.22696f
C75 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_91 VGND 1.22762f
C76 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_90 VGND 1.22562f
C77 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_89 VGND 1.22562f
C78 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_88 VGND 1.22562f
C79 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_87 VGND 1.22696f
C80 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_86 VGND 1.22562f
C81 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_85 VGND 1.22562f
C82 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_84 VGND 1.22562f
C83 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_83 VGND 1.22629f
C84 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_82 VGND 1.22696f
C85 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_81 VGND 1.22762f
C86 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_80 VGND 1.22562f
C87 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_79 VGND 1.22562f
C88 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_78 VGND 1.22629f
C89 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_77 VGND 1.22696f
C90 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_76 VGND 1.22562f
C91 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_75 VGND 1.22562f
C92 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_74 VGND 1.22562f
C93 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_73 VGND 1.22629f
C94 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_72 VGND 1.22696f
C95 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_71 VGND 1.22562f
C96 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_70 VGND 1.22562f
C97 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_69 VGND 1.22562f
C98 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_68 VGND 1.22629f
C99 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_67 VGND 1.22696f
C100 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_66 VGND 1.22762f
C101 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_65 VGND 1.22562f
C102 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_64 VGND 1.22562f
C103 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_63 VGND 1.22629f
C104 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_62 VGND 1.22696f
C105 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_61 VGND 1.22762f
C106 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_60 VGND 1.22562f
C107 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_59 VGND 1.22562f
C108 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_58 VGND 1.22629f
C109 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_57 VGND 1.22562f
C110 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_56 VGND 1.22762f
C111 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_55 VGND 1.22562f
C112 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_54 VGND 1.22562f
C113 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_53 VGND 1.22629f
C114 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_52 VGND 1.22696f
C115 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_51 VGND 1.22762f
C116 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_50 VGND 1.22562f
C117 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_49 VGND 1.22562f
C118 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_48 VGND 1.22629f
C119 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_47 VGND 1.22696f
C120 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_46 VGND 1.22562f
C121 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_45 VGND 1.22562f
C122 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_44 VGND 1.22562f
C123 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_43 VGND 1.22629f
C124 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_42 VGND 1.22696f
C125 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_41 VGND 1.22762f
C126 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_40 VGND 1.22562f
C127 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_39 VGND 1.22562f
C128 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_38 VGND 1.22629f
C129 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_37 VGND 1.22696f
C130 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2n VGND 56.048f
C131 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_35 VGND 1.22829f
C132 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_34 VGND 1.22562f
C133 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_33 VGND 1.22629f
C134 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_32 VGND 1.22696f
C135 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_31 VGND 1.22762f
C136 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_30 VGND 1.22562f
C137 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_29 VGND 1.22562f
C138 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_28 VGND 1.22629f
C139 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_27 VGND 1.22696f
C140 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_26 VGND 1.22562f
C141 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_25 VGND 1.22562f
C142 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_24 VGND 1.22562f
C143 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_23 VGND 1.22629f
C144 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_22 VGND 1.22696f
C145 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_21 VGND 1.22762f
C146 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_20 VGND 1.22562f
C147 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_19 VGND 1.22562f
C148 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_18 VGND 1.22629f
C149 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1n VGND 78.81621f
C150 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_16 VGND 1.22562f
C151 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_15 VGND 1.22562f
C152 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_14 VGND 1.22562f
C153 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_13 VGND 1.22629f
C154 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_12 VGND 1.22562f
C155 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_11 VGND 1.22762f
C156 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_10 VGND 1.22562f
C157 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_9 VGND 1.22562f
C158 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_8 VGND 1.22629f
C159 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_7 VGND 1.22696f
C160 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_6 VGND 1.22562f
C161 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_5 VGND 1.22562f
C162 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_4 VGND 1.22562f
C163 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_3 VGND 1.22629f
C164 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_2 VGND 1.22896f
C165 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_1 VGND 1.22562f
C166 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_0 VGND 1.22562f
C167 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VGND 14.3155f
C168 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VGND 4.48926f
C169 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VGND 7.66312f
C170 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VGND 7.89561f
C171 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin VGND 2.82434f
C172 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C173 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C174 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VGND 2.49069f
C175 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C176 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C177 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C178 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C179 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C180 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VGND 2.49069f
C181 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C182 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C183 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VGND 11.5086f
C184 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VGND 4.48926f
C185 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VGND 2.83622f
C186 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C187 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C188 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VGND 5.82216f
C189 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C190 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND 51.5669f
C191 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C192 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C193 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutp VGND 71.3916f
C194 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C195 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C196 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VGND 5.82216f
C197 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C198 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 VGND 33.3927f
C199 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND 75.0436f
C200 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C201 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VGND 37.237f
C202 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VGND 14.3155f
C203 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VGND 4.48926f
C204 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VGND 7.66312f
C205 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VGND 7.89561f
C206 iq_modulator_0.iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin VGND 2.82434f
C207 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.voutn VGND 77.9315f
C208 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_136 VGND 1.22562f
C209 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_135 VGND 1.22562f
C210 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_134 VGND 1.22562f
C211 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_133 VGND 1.22562f
C212 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_132 VGND 1.22696f
C213 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_131 VGND 1.22562f
C214 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_130 VGND 1.22562f
C215 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_129 VGND 1.22562f
C216 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_128 VGND 1.22629f
C217 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_127 VGND 1.22562f
C218 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_126 VGND 1.22562f
C219 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_125 VGND 1.22562f
C220 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_124 VGND 1.22562f
C221 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_123 VGND 1.22629f
C222 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_122 VGND 1.22696f
C223 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_121 VGND 1.22562f
C224 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_120 VGND 1.22562f
C225 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_119 VGND 1.22629f
C226 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_118 VGND 1.22629f
C227 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_117 VGND 1.22562f
C228 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_116 VGND 1.22562f
C229 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_115 VGND 1.22562f
C230 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_114 VGND 1.22562f
C231 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_113 VGND 1.22562f
C232 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_112 VGND 1.22696f
C233 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_111 VGND 1.22562f
C234 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_110 VGND 1.22562f
C235 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_109 VGND 1.22562f
C236 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_108 VGND 1.22629f
C237 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_107 VGND 1.22696f
C238 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_106 VGND 1.22562f
C239 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_105 VGND 1.22562f
C240 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_104 VGND 1.22562f
C241 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_103 VGND 1.22629f
C242 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_102 VGND 1.22696f
C243 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_101 VGND 1.22562f
C244 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_100 VGND 1.22562f
C245 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 VGND 39.0581f
C246 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_98 VGND 1.22629f
C247 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_97 VGND 1.22562f
C248 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_96 VGND 1.22562f
C249 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_95 VGND 1.22562f
C250 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_94 VGND 1.22562f
C251 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_93 VGND 1.22629f
C252 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_92 VGND 1.22696f
C253 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_91 VGND 1.22562f
C254 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_90 VGND 1.22562f
C255 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_89 VGND 1.22629f
C256 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_88 VGND 1.22629f
C257 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_87 VGND 1.22562f
C258 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_86 VGND 1.22562f
C259 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_85 VGND 1.22562f
C260 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_84 VGND 1.22562f
C261 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_83 VGND 1.22629f
C262 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_82 VGND 1.22696f
C263 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_81 VGND 1.22562f
C264 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_80 VGND 1.22562f
C265 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_79 VGND 1.22562f
C266 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_78 VGND 1.22629f
C267 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_77 VGND 1.22562f
C268 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_76 VGND 1.22562f
C269 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_75 VGND 1.22562f
C270 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_74 VGND 1.22562f
C271 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_73 VGND 1.22629f
C272 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_72 VGND 1.22562f
C273 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_71 VGND 1.22562f
C274 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_70 VGND 1.22562f
C275 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_69 VGND 1.22562f
C276 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_68 VGND 1.22629f
C277 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_67 VGND 1.22696f
C278 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_66 VGND 1.22562f
C279 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_65 VGND 1.22562f
C280 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_64 VGND 1.22562f
C281 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_63 VGND 1.22629f
C282 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_62 VGND 1.22696f
C283 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_61 VGND 1.22562f
C284 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_60 VGND 1.22562f
C285 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_59 VGND 1.22562f
C286 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_58 VGND 1.22562f
C287 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_57 VGND 1.22696f
C288 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_56 VGND 1.22562f
C289 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_55 VGND 1.22562f
C290 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_54 VGND 1.22562f
C291 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_53 VGND 1.22629f
C292 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_52 VGND 1.22696f
C293 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_51 VGND 1.22562f
C294 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_50 VGND 1.22562f
C295 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_49 VGND 1.22562f
C296 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_48 VGND 1.22629f
C297 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_47 VGND 1.22562f
C298 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_46 VGND 1.22562f
C299 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_45 VGND 1.22562f
C300 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_44 VGND 1.22562f
C301 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_43 VGND 1.22629f
C302 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_42 VGND 1.22696f
C303 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_41 VGND 1.22562f
C304 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_40 VGND 1.22562f
C305 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_39 VGND 1.22562f
C306 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_38 VGND 1.22629f
C307 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_37 VGND 1.22562f
C308 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC2p VGND 59.6624f
C309 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_35 VGND 1.22562f
C310 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_34 VGND 1.22562f
C311 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_33 VGND 1.22629f
C312 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_32 VGND 1.22696f
C313 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_31 VGND 1.22562f
C314 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_30 VGND 1.22562f
C315 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_29 VGND 1.22562f
C316 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_28 VGND 1.22629f
C317 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_27 VGND 1.22562f
C318 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_26 VGND 1.22562f
C319 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_25 VGND 1.22562f
C320 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_24 VGND 1.22562f
C321 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_23 VGND 1.22629f
C322 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_22 VGND 1.22696f
C323 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_21 VGND 1.22562f
C324 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_20 VGND 1.22562f
C325 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_19 VGND 1.22562f
C326 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_18 VGND 1.22629f
C327 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.vC1p VGND 80.2351f
C328 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_16 VGND 1.22562f
C329 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_15 VGND 1.22562f
C330 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_14 VGND 1.22562f
C331 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_13 VGND 1.22562f
C332 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_12 VGND 1.22696f
C333 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_11 VGND 1.22562f
C334 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_10 VGND 1.22562f
C335 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_9 VGND 1.22562f
C336 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_8 VGND 1.22629f
C337 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_7 VGND 1.22562f
C338 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_6 VGND 1.22562f
C339 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_5 VGND 1.22562f
C340 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_4 VGND 1.22562f
C341 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_3 VGND 1.22896f
C342 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_2 VGND 1.22562f
C343 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_1 VGND 1.22562f
C344 iq_modulator_0.iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_0 VGND 1.22562f
C345 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VGND 11.5065f
C346 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VGND 4.48926f
C347 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VGND 2.83622f
C348 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_136 VGND 1.22562f
C349 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_135 VGND 1.22562f
C350 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_134 VGND 1.22562f
C351 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_133 VGND 1.22629f
C352 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_132 VGND 1.22562f
C353 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_131 VGND 1.22762f
C354 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_130 VGND 1.22562f
C355 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_129 VGND 1.22562f
C356 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_128 VGND 1.22629f
C357 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_127 VGND 1.22696f
C358 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_126 VGND 1.22562f
C359 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_125 VGND 1.22562f
C360 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_124 VGND 1.22562f
C361 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_123 VGND 1.22629f
C362 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_122 VGND 1.22696f
C363 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_121 VGND 1.22762f
C364 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_120 VGND 1.22562f
C365 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_119 VGND 1.22562f
C366 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_118 VGND 1.22562f
C367 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_117 VGND 1.22696f
C368 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_116 VGND 1.22562f
C369 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_115 VGND 1.22562f
C370 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_114 VGND 1.22562f
C371 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_113 VGND 1.22629f
C372 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_112 VGND 1.22562f
C373 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_111 VGND 1.22762f
C374 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_110 VGND 1.22562f
C375 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_109 VGND 1.22562f
C376 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_108 VGND 1.22629f
C377 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_107 VGND 1.22696f
C378 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_106 VGND 1.22762f
C379 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_105 VGND 1.22562f
C380 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_104 VGND 1.22562f
C381 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_103 VGND 1.22629f
C382 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_102 VGND 1.22696f
C383 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_101 VGND 1.22762f
C384 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_100 VGND 1.22562f
C385 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_98 VGND 1.22629f
C386 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_97 VGND 1.22696f
C387 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_96 VGND 1.22562f
C388 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_95 VGND 1.22562f
C389 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_94 VGND 1.22562f
C390 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_93 VGND 1.22629f
C391 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_92 VGND 1.22696f
C392 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_91 VGND 1.22762f
C393 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_90 VGND 1.22562f
C394 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_89 VGND 1.22562f
C395 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_88 VGND 1.22562f
C396 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_87 VGND 1.22696f
C397 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_86 VGND 1.22562f
C398 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_85 VGND 1.22562f
C399 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_84 VGND 1.22562f
C400 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_83 VGND 1.22629f
C401 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_82 VGND 1.22696f
C402 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_81 VGND 1.22762f
C403 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_80 VGND 1.22562f
C404 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_79 VGND 1.22562f
C405 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_78 VGND 1.22629f
C406 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_77 VGND 1.22696f
C407 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_76 VGND 1.22562f
C408 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_75 VGND 1.22562f
C409 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_74 VGND 1.22562f
C410 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_73 VGND 1.22629f
C411 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_72 VGND 1.22696f
C412 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_71 VGND 1.22562f
C413 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_70 VGND 1.22562f
C414 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_69 VGND 1.22562f
C415 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_68 VGND 1.22629f
C416 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_67 VGND 1.22696f
C417 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_66 VGND 1.22762f
C418 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_65 VGND 1.22562f
C419 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_64 VGND 1.22562f
C420 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_63 VGND 1.22629f
C421 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_62 VGND 1.22696f
C422 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_61 VGND 1.22762f
C423 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_60 VGND 1.22562f
C424 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_59 VGND 1.22562f
C425 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_58 VGND 1.22629f
C426 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_57 VGND 1.22562f
C427 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_56 VGND 1.22762f
C428 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_55 VGND 1.22562f
C429 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_54 VGND 1.22562f
C430 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_53 VGND 1.22629f
C431 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_52 VGND 1.22696f
C432 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_51 VGND 1.22762f
C433 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_50 VGND 1.22562f
C434 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_49 VGND 1.22562f
C435 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_48 VGND 1.22629f
C436 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_47 VGND 1.22696f
C437 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_46 VGND 1.22562f
C438 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_45 VGND 1.22562f
C439 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_44 VGND 1.22562f
C440 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_43 VGND 1.22629f
C441 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_42 VGND 1.22696f
C442 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_41 VGND 1.22762f
C443 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_40 VGND 1.22562f
C444 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_39 VGND 1.22562f
C445 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_38 VGND 1.22629f
C446 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_37 VGND 1.22696f
C447 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n VGND 59.4865f
C448 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_35 VGND 1.22829f
C449 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_34 VGND 1.22562f
C450 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_33 VGND 1.22629f
C451 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_32 VGND 1.22696f
C452 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_31 VGND 1.22762f
C453 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_30 VGND 1.22562f
C454 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_29 VGND 1.22562f
C455 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_28 VGND 1.22629f
C456 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_27 VGND 1.22696f
C457 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_26 VGND 1.22562f
C458 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_25 VGND 1.22562f
C459 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_24 VGND 1.22562f
C460 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_23 VGND 1.22629f
C461 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_22 VGND 1.22696f
C462 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_21 VGND 1.22762f
C463 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_20 VGND 1.22562f
C464 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_19 VGND 1.22562f
C465 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_18 VGND 1.22629f
C466 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n VGND 79.4888f
C467 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_16 VGND 1.22562f
C468 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_15 VGND 1.22562f
C469 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_14 VGND 1.22562f
C470 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_13 VGND 1.22629f
C471 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_12 VGND 1.22562f
C472 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_11 VGND 1.22762f
C473 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_10 VGND 1.22562f
C474 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_9 VGND 1.22562f
C475 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_8 VGND 1.22629f
C476 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_7 VGND 1.22696f
C477 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_6 VGND 1.22562f
C478 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_5 VGND 1.22562f
C479 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_4 VGND 1.22562f
C480 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_3 VGND 1.22629f
C481 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_2 VGND 1.22896f
C482 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_1 VGND 1.22562f
C483 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_0 VGND 1.22562f
C484 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VGND 14.3155f
C485 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VGND 4.48926f
C486 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VGND 7.66312f
C487 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VGND 7.89561f
C488 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin VGND 2.82434f
C489 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C490 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C491 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VGND 2.49069f
C492 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C493 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C494 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C495 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C496 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C497 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VGND 2.49069f
C498 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C499 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VGND 3.36642f
C500 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VGND 11.5086f
C501 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VGND 4.48926f
C502 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VGND 2.83622f
C503 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C504 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C505 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VGND 5.82216f
C506 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C507 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VGND 51.5669f
C508 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C509 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C510 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VGND 74.2324f
C511 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C512 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C513 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VGND 5.82216f
C514 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C515 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 VGND 36.4777f
C516 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VGND 75.0436f
C517 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VGND 7.84314f
C518 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VGND 37.237f
C519 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VGND 14.3155f
C520 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VGND 4.48926f
C521 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VGND 7.66312f
C522 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VGND 7.89561f
C523 iq_modulator_0.iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin VGND 2.82434f
C524 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VGND 74.9539f
C525 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_136 VGND 1.22562f
C526 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_135 VGND 1.22562f
C527 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_134 VGND 1.22562f
C528 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_133 VGND 1.22562f
C529 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_132 VGND 1.22696f
C530 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_131 VGND 1.22562f
C531 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_130 VGND 1.22562f
C532 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_129 VGND 1.22562f
C533 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_128 VGND 1.22629f
C534 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_127 VGND 1.22562f
C535 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_126 VGND 1.22562f
C536 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_125 VGND 1.22562f
C537 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_124 VGND 1.22562f
C538 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_123 VGND 1.22629f
C539 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_122 VGND 1.22696f
C540 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_121 VGND 1.22562f
C541 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_120 VGND 1.22562f
C542 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_119 VGND 1.22629f
C543 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_118 VGND 1.22629f
C544 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_117 VGND 1.22562f
C545 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_116 VGND 1.22562f
C546 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_115 VGND 1.22562f
C547 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_114 VGND 1.22562f
C548 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_113 VGND 1.22562f
C549 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_112 VGND 1.22696f
C550 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_111 VGND 1.22562f
C551 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_110 VGND 1.22562f
C552 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_109 VGND 1.22562f
C553 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_108 VGND 1.22629f
C554 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_107 VGND 1.22696f
C555 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_106 VGND 1.22562f
C556 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_105 VGND 1.22562f
C557 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_104 VGND 1.22562f
C558 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_103 VGND 1.22629f
C559 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_102 VGND 1.22696f
C560 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_101 VGND 1.22562f
C561 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_100 VGND 1.22562f
C562 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 VGND 36.1864f
C563 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_98 VGND 1.22629f
C564 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_97 VGND 1.22562f
C565 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_96 VGND 1.22562f
C566 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_95 VGND 1.22562f
C567 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_94 VGND 1.22562f
C568 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_93 VGND 1.22629f
C569 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_92 VGND 1.22696f
C570 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_91 VGND 1.22562f
C571 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_90 VGND 1.22562f
C572 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_89 VGND 1.22629f
C573 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_88 VGND 1.22629f
C574 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_87 VGND 1.22562f
C575 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_86 VGND 1.22562f
C576 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_85 VGND 1.22562f
C577 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_84 VGND 1.22562f
C578 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_83 VGND 1.22629f
C579 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_82 VGND 1.22696f
C580 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_81 VGND 1.22562f
C581 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_80 VGND 1.22562f
C582 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_79 VGND 1.22562f
C583 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_78 VGND 1.22629f
C584 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_77 VGND 1.22562f
C585 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_76 VGND 1.22562f
C586 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_75 VGND 1.22562f
C587 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_74 VGND 1.22562f
C588 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_73 VGND 1.22629f
C589 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_72 VGND 1.22562f
C590 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_71 VGND 1.22562f
C591 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_70 VGND 1.22562f
C592 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_69 VGND 1.22562f
C593 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_68 VGND 1.22629f
C594 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_67 VGND 1.22696f
C595 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_66 VGND 1.22562f
C596 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_65 VGND 1.22562f
C597 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_64 VGND 1.22562f
C598 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_63 VGND 1.22629f
C599 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_62 VGND 1.22696f
C600 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_61 VGND 1.22562f
C601 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_60 VGND 1.22562f
C602 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_59 VGND 1.22562f
C603 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_58 VGND 1.22562f
C604 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_57 VGND 1.22696f
C605 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_56 VGND 1.22562f
C606 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_55 VGND 1.22562f
C607 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_54 VGND 1.22562f
C608 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_53 VGND 1.22629f
C609 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_52 VGND 1.22696f
C610 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_51 VGND 1.22562f
C611 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_50 VGND 1.22562f
C612 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_49 VGND 1.22562f
C613 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_48 VGND 1.22629f
C614 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_47 VGND 1.22562f
C615 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_46 VGND 1.22562f
C616 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_45 VGND 1.22562f
C617 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_44 VGND 1.22562f
C618 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_43 VGND 1.22629f
C619 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_42 VGND 1.22696f
C620 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_41 VGND 1.22562f
C621 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_40 VGND 1.22562f
C622 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_39 VGND 1.22562f
C623 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_38 VGND 1.22629f
C624 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_37 VGND 1.22562f
C625 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p VGND 56.026f
C626 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_35 VGND 1.22562f
C627 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_34 VGND 1.22562f
C628 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_33 VGND 1.22629f
C629 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_32 VGND 1.22696f
C630 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_31 VGND 1.22562f
C631 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_30 VGND 1.22562f
C632 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_29 VGND 1.22562f
C633 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_28 VGND 1.22629f
C634 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_27 VGND 1.22562f
C635 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_26 VGND 1.22562f
C636 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_25 VGND 1.22562f
C637 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_24 VGND 1.22562f
C638 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_23 VGND 1.22629f
C639 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_22 VGND 1.22696f
C640 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_21 VGND 1.22562f
C641 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_20 VGND 1.22562f
C642 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_19 VGND 1.22562f
C643 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_18 VGND 1.22629f
C644 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p VGND 78.8372f
C645 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_16 VGND 1.22562f
C646 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_15 VGND 1.22562f
C647 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_14 VGND 1.22562f
C648 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_13 VGND 1.22562f
C649 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_12 VGND 1.22696f
C650 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_11 VGND 1.22562f
C651 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_10 VGND 1.22562f
C652 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_9 VGND 1.22562f
C653 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_8 VGND 1.22629f
C654 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_7 VGND 1.22562f
C655 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_6 VGND 1.22562f
C656 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_5 VGND 1.22562f
C657 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_4 VGND 1.22562f
C658 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_3 VGND 1.22896f
C659 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_2 VGND 1.22562f
C660 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_1 VGND 1.22562f
C661 iq_modulator_0.iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_0 VGND 1.22562f
.ends

