magic
tech sky130A
magscale 1 2
timestamp 1762641840
<< locali >>
rect 4990 2730 8250 3940
rect 5325 2630 8250 2730
rect 5325 2625 5355 2630
rect 5325 820 8250 925
rect 4990 30 8250 820
rect 4990 -1440 8250 -230
rect 5325 -1610 8250 -1440
rect 5325 -3250 5685 -3245
rect 5325 -3355 8250 -3250
rect 4990 -4140 8250 -3355
<< metal1 >>
rect 2130 3760 2705 3970
rect 4935 3925 7280 3940
rect 4935 3700 6675 3925
rect 4990 3685 6675 3700
rect 7265 3685 7280 3925
rect 4990 3670 7280 3685
rect 0 1775 120 1865
rect 4990 285 6290 300
rect 4990 270 5685 285
rect 4935 45 5685 270
rect 6275 45 6290 285
rect 4935 30 6290 45
rect 4935 -245 7280 -230
rect 4935 -470 6675 -245
rect 4990 -485 6675 -470
rect 7265 -485 7280 -245
rect 4990 -500 7280 -485
rect 0 -2410 120 -2285
rect 4990 -3885 6755 -3870
rect 4990 -3900 6150 -3885
rect 2265 -4140 2550 -4030
rect 4935 -4125 6150 -3900
rect 6740 -4125 6755 -3885
rect 4935 -4140 6755 -4125
<< via1 >>
rect 6675 3685 7265 3925
rect 5335 2460 8240 2515
rect 5515 1515 5730 1625
rect 5685 45 6275 285
rect 6675 -485 7265 -245
rect 5335 -1710 8240 -1655
rect 5515 -2660 5675 -2550
rect 6150 -4125 6740 -3885
<< metal2 >>
rect 6660 3925 7280 3940
rect 6660 3685 6675 3925
rect 7265 3685 7280 3925
rect 6660 3670 7280 3685
rect 5080 2570 5200 2765
rect 5080 2515 8250 2570
rect 5080 2460 5335 2515
rect 8240 2460 8250 2515
rect 5080 2450 8250 2460
rect 5080 1625 5740 1635
rect 5080 1515 5515 1625
rect 5730 1515 5740 1625
rect 5080 1505 5740 1515
rect 5080 785 5200 1505
rect 5670 285 6290 300
rect 5670 45 5685 285
rect 6275 45 6290 285
rect 5670 30 6290 45
rect 6660 -245 7280 -230
rect 6660 -485 6675 -245
rect 7265 -485 7280 -245
rect 6660 -500 7280 -485
rect 5080 -1600 5200 -1405
rect 5080 -1655 8250 -1600
rect 5080 -1710 5335 -1655
rect 8240 -1710 8250 -1655
rect 5080 -1720 8250 -1710
rect 5025 -2550 5685 -2540
rect 5025 -2660 5515 -2550
rect 5675 -2660 5685 -2550
rect 5025 -2670 5685 -2660
rect 5025 -3385 5145 -2670
rect 6135 -3885 6755 -3870
rect 6135 -4125 6150 -3885
rect 6740 -4125 6755 -3885
rect 6135 -4140 6755 -4125
<< via2 >>
rect 6675 3685 7265 3925
rect 5685 45 6275 285
rect 6675 -485 7265 -245
rect 6150 -4125 6740 -3885
<< metal3 >>
rect 875 -3970 1185 2470
rect 1795 -3080 2105 3550
rect 3635 -3970 3945 2470
rect 4990 2390 5810 3995
rect 6660 3925 7280 3940
rect 6660 3685 6675 3925
rect 7265 3685 7280 3925
rect 4990 1120 5300 2390
rect 5670 285 6290 300
rect 5670 45 5685 285
rect 6275 45 6290 285
rect 5670 -840 6290 45
rect 6660 -245 7280 3685
rect 6660 -485 6675 -245
rect 7265 -485 7280 -245
rect 6660 -500 7280 -485
rect 5670 -1460 6755 -840
rect 4990 -3045 5300 -1775
rect 4990 -4195 5810 -3045
rect 6135 -3885 6755 -1460
rect 7670 -3050 9030 2395
rect 6135 -4125 6150 -3885
rect 6740 -4125 6755 -3885
rect 6135 -4140 6755 -4125
use lo_logic  lo_logic_0 lo_logic
timestamp 1762641840
transform 1 0 195 0 1 2060
box -195 -2030 5005 1880
use lo_logic  lo_logic_1
timestamp 1762641840
transform 1 0 195 0 1 -2110
box -195 -2030 5005 1880
use transmission_gate_w_dummy  transmission_gate_w_dummy_0 transmission_gate_w_dummy
timestamp 1762641840
transform 1 0 5340 0 1 1640
box -40 -720 2935 990
use transmission_gate_w_dummy  transmission_gate_w_dummy_2
timestamp 1762641840
transform 1 0 5340 0 1 -2530
box -40 -720 2935 990
<< labels >>
flabel metal1 2405 3865 2405 3865 0 FreeSans 1600 0 0 0 VDD
port 9 nsew
flabel metal3 8800 -235 8800 -235 0 FreeSans 800 0 0 0 vout_RF
port 19 nsew
flabel metal1 2400 -4085 2400 -4085 0 FreeSans 1600 0 0 0 VSS
port 21 nsew
flabel metal1 55 1825 55 1825 0 FreeSans 800 0 0 0 vinn_LO
port 76 nsew
flabel metal1 55 -2355 55 -2355 0 FreeSans 800 0 0 0 vinp_LO
port 78 nsew
flabel metal3 5385 3965 5385 3965 0 FreeSans 800 0 0 0 vinn_IF
port 80 nsew
flabel metal3 5375 -4165 5375 -4165 0 FreeSans 800 0 0 0 vinp_IF
port 82 nsew
<< end >>
