* PEX produced on Fri Nov  7 02:57:23 PM CET 2025 using /foss/tools/sak/iic-pex.sh with m=1 and s=1
* NGSPICE file created from third_order_mfb_lp_filter_wo_C.ext - technology: sky130A

.subckt third_order_mfb_lp_filter_wo_C_pex vinp vinn vC1p vC1n vC2n vC2p di_filter_ota_en
+ voutn voutp VDD VSS
X0 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_61 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_62 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_2 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_3 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X2 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_111 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_110 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X3 ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X4 voutp resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X5 ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X6 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_15 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_14 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X7 VDD ota_core_hybrid_bm_0.ota_core_en_n ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X8 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_77 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_76 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X9 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X10 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_128 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_127 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X11 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_125 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_126 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X12 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X13 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_78 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_79 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X14 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_68 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_69 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X15 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 voutp ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X16 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_26 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_25 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X17 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_29 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_30 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X18 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_67 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_68 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X19 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_21 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_22 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X20 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout voutp ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X21 ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 voutp VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X22 ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout voutn VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X23 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_108 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_109 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X24 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_50 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_49 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X25 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_21 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_20 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X26 VDD ota_core_hybrid_bm_0.ota_core_en_n ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X27 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_83 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_82 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X28 ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout voutp VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X29 ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 voutn ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X30 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_38 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_39 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X31 ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X32 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_35 vC2n VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X33 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_117 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_116 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X34 voutp ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X35 ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X36 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_73 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_74 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X37 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_27 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_28 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X38 ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 voutn VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X39 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_122 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_121 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X40 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_3 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_4 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X41 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_72 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_73 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X42 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_62 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_63 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X43 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_104 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_105 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X44 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_20 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_19 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X45 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout voutp ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X46 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X47 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_89 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_88 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X48 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_131 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_132 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X49 ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X50 voutn resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X51 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_64 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_63 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X52 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_123 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_122 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X53 ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X54 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_54 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_53 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X55 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X56 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_134 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_135 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X57 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_96 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_95 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X58 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_33 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_34 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X59 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_10 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_11 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X60 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_86 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_85 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X61 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_0 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_1 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X62 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_42 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_43 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X63 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_27 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_26 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X64 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_32 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_33 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X65 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 voutp ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X66 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_66 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_67 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X67 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_126 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_125 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X68 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_105 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_106 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X69 voutn ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X70 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_41 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_42 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X71 ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X72 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_116 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_115 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X73 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_56 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_57 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X74 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_34 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_33 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X75 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_79 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_80 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X76 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X77 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_129 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_128 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X78 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_24 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_23 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X79 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_71 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_72 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X80 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_9 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_10 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X81 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_47 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_48 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X82 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout voutp ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X83 ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 voutp VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X84 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_33 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_32 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X85 VSS VDD ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X86 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_25 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_24 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X87 ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout voutp VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X88 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_58 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_57 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X89 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_95 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_94 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X90 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_48 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_47 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X91 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_1 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_0 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X92 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_90 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_89 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X93 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_4 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_5 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X94 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_80 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_79 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X95 vC2p resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_37 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X96 ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X97 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_26 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_27 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X98 voutn ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X99 voutp ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X100 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_85 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_86 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X101 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_39 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_40 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X102 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_77 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_78 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X103 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_15 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_16 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X104 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout voutn ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X105 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_53 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_54 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X106 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_120 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_119 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X107 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_45 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_46 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X108 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_39 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_38 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X109 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout voutp ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X110 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_70 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_71 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X111 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_110 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_109 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X112 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_101 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_100 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X113 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_31 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_30 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X114 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_28 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_27 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X115 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_102 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_103 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X116 ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X117 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_18 vC1p VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X118 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_111 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_112 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X119 ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X120 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_135 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_134 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X121 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X122 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_52 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_51 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X123 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_83 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_84 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X124 ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X125 VSS VDD ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X126 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_132 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_133 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X127 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_94 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_93 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X128 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X129 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_40 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_41 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X130 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_7 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_6 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X131 voutn ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X132 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_117 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_118 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X133 ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X134 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_91 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_92 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X135 VSS VDD ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X136 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X137 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_124 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_123 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X138 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_64 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_65 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X139 VSS VDD ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X140 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_22 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_21 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X141 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_96 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_97 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X142 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_59 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_60 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X143 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_12 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_11 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X144 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_109 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_108 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X145 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_45 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_44 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X146 VDD ota_core_hybrid_bm_0.ota_core_en_n ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X147 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_51 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_52 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X148 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X149 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_37 vC2n VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X150 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_75 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_74 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X151 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_13 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_12 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X152 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_51 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_50 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X153 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_5 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_4 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X154 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_136 voutn VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X155 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_123 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_124 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X156 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_88 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_87 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X157 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_126 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_127 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X158 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_97 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_98 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X159 voutn ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X160 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_34 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_35 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X161 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_89 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_90 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X162 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout voutn ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X163 ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X164 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_65 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_66 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X165 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout voutp ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X166 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_57 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_58 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X167 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_43 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_42 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X168 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_81 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_80 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X169 ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X170 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_118 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_117 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X171 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_19 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_18 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X172 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_11 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_10 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X173 ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X174 ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X175 ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X176 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_100 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_101 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X177 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_49 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_48 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X178 VSS VDD ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X179 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_16 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_15 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X180 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X181 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_103 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_104 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X182 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_95 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_96 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X183 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X184 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_115 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_114 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X185 VDD ota_core_hybrid_bm_0.ota_core_en_n ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X186 ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X187 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X188 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X189 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_63 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_64 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X190 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_82 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_81 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X191 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_57 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_56 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X192 ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X193 VSS VDD ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X194 ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 voutn VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X195 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_129 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_130 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X196 VDD ota_core_hybrid_bm_0.ota_core_en_n ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X197 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_98 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X198 VDD ota_core_hybrid_bm_0.ota_core_en_n ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X199 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_14 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_13 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X200 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_1 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_2 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X201 voutn resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X202 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_112 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_111 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X203 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_121 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_120 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X204 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X205 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_94 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_95 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X206 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_10 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_9 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X207 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_87 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_86 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X208 ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 voutn ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X209 ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X210 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_42 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_41 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X211 ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 voutn VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X212 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_63 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_62 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X213 vC1n resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_16 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X214 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_128 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_129 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X215 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_55 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_54 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X216 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_135 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_136 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X217 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_101 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_102 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X218 ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X219 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_7 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_8 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X220 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout voutp ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X221 VSS VDD ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X222 ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout voutn VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X223 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_69 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_70 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X224 voutn resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X225 ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X226 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_60 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_61 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X227 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_50 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_51 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X228 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_93 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_92 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X229 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_92 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_93 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X230 ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X231 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_8 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_7 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X232 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_69 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_68 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X233 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_23 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_22 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X234 ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X235 VDD ota_core_hybrid_bm_0.ota_core_en_n ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X236 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_61 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_60 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X237 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X238 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X239 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_127 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_126 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X240 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_13 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_14 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X241 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_122 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_123 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X242 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_84 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_83 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X243 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_75 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_76 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X244 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X245 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_74 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_73 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X246 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_30 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_31 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X247 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X248 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_98 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X249 ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X250 VDD ota_core_hybrid_bm_0.ota_core_en_n ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X251 ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 voutn VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X252 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_20 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_21 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X253 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_29 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_28 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X254 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_54 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_55 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X255 VSS VDD ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X256 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_114 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_113 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X257 ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 voutp VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X258 VSS di_filter_ota_en ota_core_hybrid_bm_0.ota_core_en_n VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X259 voutn resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X260 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_86 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_87 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X261 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_133 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_132 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X262 VSS VDD ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X263 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_2 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_1 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X264 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_125 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_124 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X265 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_44 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_43 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X266 ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 voutn ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X267 ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X268 voutp resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X269 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=23.49 ps=177.66 w=3 l=1
X270 ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 voutn VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X271 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 voutp ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X272 voutp ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X273 ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X274 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_46 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_45 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X275 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_67 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_66 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X276 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_78 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_77 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X277 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_116 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_117 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X278 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_68 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_67 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X279 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_24 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_25 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X280 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_19 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_20 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X281 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X282 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X283 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_14 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_15 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X284 ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout voutn VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X285 VDD ota_core_hybrid_bm_0.ota_core_en_n ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X286 voutn resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X287 ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X288 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_81 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_82 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X289 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X290 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_131 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_130 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X291 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_105 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_104 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X292 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_108 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_107 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X293 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_35 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_34 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X294 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_58 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_59 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X295 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_73 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_72 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X296 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_90 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_91 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X297 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_6 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_5 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X298 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_38 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_37 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X299 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_25 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_26 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X300 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_87 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_88 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X301 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_130 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_131 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X302 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_107 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_106 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X303 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X304 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_72 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_71 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X305 ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X306 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_120 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_121 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X307 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_62 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_61 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X308 ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X309 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_41 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_40 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X310 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_28 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_29 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X311 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_121 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_122 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X312 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_104 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_103 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X313 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_79 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_78 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X314 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_18 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_19 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X315 VDD ota_core_hybrid_bm_0.ota_core_en_n ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X316 ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 voutp VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X317 VDD di_filter_ota_en ota_core_hybrid_bm_0.ota_core_en_n VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X318 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X319 VDD ota_core_hybrid_bm_0.ota_core_en_n ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X320 ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout voutn VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X321 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_52 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_53 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X322 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_93 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_94 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X323 voutp resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_136 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X324 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_84 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_85 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X325 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_113 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_112 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X326 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_0 vinp VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X327 voutp resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X328 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=70.47 ps=501.66 w=9 l=1
X329 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 voutp ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X330 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_32 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_31 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X331 ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X332 voutn ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X333 voutp ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X334 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_127 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_128 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X335 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout voutn ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X336 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_47 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_46 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X337 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_124 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_125 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X338 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X339 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_31 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_32 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X340 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_76 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_75 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X341 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X342 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_114 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_115 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X343 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_66 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_65 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X344 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X345 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_22 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_23 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X346 ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 voutn ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X347 vinn resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_0 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X348 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_98 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_97 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X349 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_12 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_13 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X350 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_119 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_118 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X351 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_44 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_45 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X352 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_85 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_84 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X353 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_133 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_134 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X354 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_106 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_105 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X355 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_46 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_47 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X356 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X357 ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout voutp VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X358 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_53 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_52 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X359 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout voutn ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X360 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X361 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_88 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_89 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X362 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_4 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_3 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X363 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_37 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_38 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X364 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0 ps=0 w=3 l=1
X365 vC2p resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_35 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X366 vC2n resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_100 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X367 ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X368 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_5 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_6 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X369 ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X370 ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X371 voutp ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X372 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_70 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_69 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X373 ota_core_hybrid_bm_0.ota_core_en_n di_filter_ota_en VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X374 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_60 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_59 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X375 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_91 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_90 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X376 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_118 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_119 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X377 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_102 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_101 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X378 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_109 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_110 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X379 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_16 vC1p VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X380 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_92 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_91 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X381 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_6 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_7 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X382 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_59 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_58 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X383 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X384 ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout voutp VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X385 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_43 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_44 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X386 ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout voutn VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X387 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 voutp ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X388 voutp resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X389 VSS di_filter_ota_en ota_core_hybrid_bm_0.ota_core_en_n VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X390 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_132 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_131 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X391 voutn ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X392 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_82 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_83 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X393 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_40 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_39 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X394 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout voutn ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X395 ota_core_hybrid_bm_0.ota_core_en_n di_filter_ota_en VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X396 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_30 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_29 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X397 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_115 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_116 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X398 ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 voutp VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X399 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X400 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_107 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_108 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X401 ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 voutn ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X402 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_11 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_12 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X403 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_112 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_113 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X404 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_49 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_50 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X405 ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X406 voutp resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X407 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_48 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_49 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X408 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_97 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_96 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X409 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_80 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_81 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X410 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_3 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_2 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X411 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X412 VSS VDD ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X413 ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout voutp VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X414 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_65 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_64 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X415 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout voutn ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X416 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X417 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_113 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_114 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X418 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X419 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X420 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=0 ps=0 w=9 l=1
X421 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_136 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_135 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X422 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_76 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_77 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X423 ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X424 vC1n resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_18 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X425 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_55 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_56 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X426 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_110 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_111 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X427 voutp ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X428 ota_core_hybrid_bm_0.ota_core_en_n di_filter_ota_en VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X429 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_103 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_102 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X430 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_9 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_8 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X431 ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout voutn VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X432 VSS VDD ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X433 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_8 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_9 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X434 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_106 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_107 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X435 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_71 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_70 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X436 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_100 vC2p VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X437 ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout voutp VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X438 ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 voutn ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X439 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 voutp ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X440 ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X441 VDD di_filter_ota_en ota_core_hybrid_bm_0.ota_core_en_n VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X442 voutp resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X443 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_134 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_133 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X444 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_23 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_24 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X445 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_74 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_75 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X446 ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 voutn VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X447 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_130 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_129 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X448 ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 voutp VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X449 ota_core_hybrid_bm_0.ota_core_en_n di_filter_ota_en VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X450 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X451 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_119 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_120 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X452 ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X453 voutn resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X454 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X455 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_56 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_55 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
C0 vC2n VSS 8.47651f
C1 vC1n VSS 1.23726f
C2 vinn VSS 3.70189f
C3 voutp VSS 43.7785f
C4 di_filter_ota_en VSS 4.83684f
C5 voutn VSS 47.1455f
C6 vC2p VSS 8.43064f
C7 vC1p VSS 1.24123f
C8 vinp VSS 3.69855f
C9 VDD VSS 0.35571p
C10 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_136 VSS 1.22562f
C11 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_135 VSS 1.22562f
C12 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_134 VSS 1.22562f
C13 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_133 VSS 1.22629f
C14 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_132 VSS 1.22562f
C15 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_131 VSS 1.22762f
C16 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_130 VSS 1.22562f
C17 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_129 VSS 1.22562f
C18 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_128 VSS 1.22629f
C19 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_127 VSS 1.22696f
C20 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_126 VSS 1.22562f
C21 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_125 VSS 1.22562f
C22 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_124 VSS 1.22562f
C23 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_123 VSS 1.22629f
C24 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_122 VSS 1.22696f
C25 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_121 VSS 1.22762f
C26 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_120 VSS 1.22562f
C27 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_119 VSS 1.22562f
C28 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_118 VSS 1.22562f
C29 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_117 VSS 1.22696f
C30 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_116 VSS 1.22562f
C31 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_115 VSS 1.22562f
C32 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_114 VSS 1.22562f
C33 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_113 VSS 1.22629f
C34 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_112 VSS 1.22562f
C35 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_111 VSS 1.22762f
C36 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_110 VSS 1.22562f
C37 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_109 VSS 1.22562f
C38 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_108 VSS 1.22629f
C39 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_107 VSS 1.22696f
C40 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_106 VSS 1.22762f
C41 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_105 VSS 1.22562f
C42 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_104 VSS 1.22562f
C43 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_103 VSS 1.22629f
C44 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_102 VSS 1.22696f
C45 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_101 VSS 1.22762f
C46 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_100 VSS 1.22562f
C47 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_98 VSS 1.22629f
C48 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_97 VSS 1.22696f
C49 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_96 VSS 1.22562f
C50 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_95 VSS 1.22562f
C51 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_94 VSS 1.22562f
C52 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_93 VSS 1.22629f
C53 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_92 VSS 1.22696f
C54 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_91 VSS 1.22762f
C55 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_90 VSS 1.22562f
C56 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_89 VSS 1.22562f
C57 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_88 VSS 1.22562f
C58 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_87 VSS 1.22696f
C59 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_86 VSS 1.22562f
C60 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_85 VSS 1.22562f
C61 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_84 VSS 1.22562f
C62 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_83 VSS 1.22629f
C63 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_82 VSS 1.22696f
C64 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_81 VSS 1.22762f
C65 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_80 VSS 1.22562f
C66 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_79 VSS 1.22562f
C67 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_78 VSS 1.22629f
C68 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_77 VSS 1.22696f
C69 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_76 VSS 1.22562f
C70 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_75 VSS 1.22562f
C71 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_74 VSS 1.22562f
C72 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_73 VSS 1.22629f
C73 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_72 VSS 1.22696f
C74 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_71 VSS 1.22562f
C75 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_70 VSS 1.22562f
C76 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_69 VSS 1.22562f
C77 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_68 VSS 1.22629f
C78 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_67 VSS 1.22696f
C79 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_66 VSS 1.22762f
C80 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_65 VSS 1.22562f
C81 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_64 VSS 1.22562f
C82 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_63 VSS 1.22629f
C83 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_62 VSS 1.22696f
C84 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_61 VSS 1.22762f
C85 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_60 VSS 1.22562f
C86 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_59 VSS 1.22562f
C87 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_58 VSS 1.22629f
C88 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_57 VSS 1.22562f
C89 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_56 VSS 1.22762f
C90 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_55 VSS 1.22562f
C91 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_54 VSS 1.22562f
C92 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_53 VSS 1.22629f
C93 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_52 VSS 1.22696f
C94 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_51 VSS 1.22762f
C95 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_50 VSS 1.22562f
C96 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_49 VSS 1.22562f
C97 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_48 VSS 1.22629f
C98 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_47 VSS 1.22696f
C99 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_46 VSS 1.22562f
C100 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_45 VSS 1.22562f
C101 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_44 VSS 1.22562f
C102 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_43 VSS 1.22629f
C103 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_42 VSS 1.22696f
C104 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_41 VSS 1.22762f
C105 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_40 VSS 1.22562f
C106 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_39 VSS 1.22562f
C107 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_38 VSS 1.22629f
C108 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_37 VSS 1.22696f
C109 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_35 VSS 1.22829f
C110 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_34 VSS 1.22562f
C111 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_33 VSS 1.22629f
C112 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_32 VSS 1.22696f
C113 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_31 VSS 1.22762f
C114 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_30 VSS 1.22562f
C115 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_29 VSS 1.22562f
C116 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_28 VSS 1.22629f
C117 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_27 VSS 1.22696f
C118 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_26 VSS 1.22562f
C119 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_25 VSS 1.22562f
C120 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_24 VSS 1.22562f
C121 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_23 VSS 1.22629f
C122 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_22 VSS 1.22696f
C123 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_21 VSS 1.22762f
C124 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_20 VSS 1.22562f
C125 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_19 VSS 1.22562f
C126 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_18 VSS 1.22629f
C127 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_16 VSS 1.22562f
C128 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_15 VSS 1.22562f
C129 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_14 VSS 1.22562f
C130 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_13 VSS 1.22629f
C131 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_12 VSS 1.22562f
C132 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_11 VSS 1.22762f
C133 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_10 VSS 1.22562f
C134 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_9 VSS 1.22562f
C135 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_8 VSS 1.22629f
C136 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_7 VSS 1.22696f
C137 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_6 VSS 1.22562f
C138 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_5 VSS 1.22562f
C139 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_4 VSS 1.22562f
C140 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_3 VSS 1.22629f
C141 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_2 VSS 1.22896f
C142 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_1 VSS 1.22562f
C143 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_0 VSS 1.22562f
C144 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS 3.36642f
C145 ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS 3.36642f
C146 ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VSS 2.49069f
C147 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS 3.36642f
C148 ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS 3.36642f
C149 ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS 3.36642f
C150 ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS 3.36642f
C151 ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS 3.36642f
C152 ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VSS 2.49069f
C153 ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS 3.36642f
C154 ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS 3.36642f
C155 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VSS 7.84314f
C156 ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VSS 7.84314f
C157 ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VSS 5.82216f
C158 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VSS 7.84314f
C159 ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VSS 51.5669f
C160 ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VSS 7.84314f
C161 ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VSS 7.84314f
C162 ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VSS 7.84314f
C163 ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VSS 7.84314f
C164 ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VSS 5.82216f
C165 ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VSS 7.84314f
C166 resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 VSS 25.9659f
C167 ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS 75.0436f
C168 ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VSS 7.84314f
C169 ota_core_hybrid_bm_0.ota_core_en_n VSS 37.237f
C170 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_136 VSS 1.22562f
C171 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_135 VSS 1.22562f
C172 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_134 VSS 1.22562f
C173 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_133 VSS 1.22562f
C174 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_132 VSS 1.22696f
C175 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_131 VSS 1.22562f
C176 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_130 VSS 1.22562f
C177 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_129 VSS 1.22562f
C178 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_128 VSS 1.22629f
C179 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_127 VSS 1.22562f
C180 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_126 VSS 1.22562f
C181 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_125 VSS 1.22562f
C182 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_124 VSS 1.22562f
C183 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_123 VSS 1.22629f
C184 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_122 VSS 1.22696f
C185 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_121 VSS 1.22562f
C186 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_120 VSS 1.22562f
C187 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_119 VSS 1.22629f
C188 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_118 VSS 1.22629f
C189 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_117 VSS 1.22562f
C190 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_116 VSS 1.22562f
C191 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_115 VSS 1.22562f
C192 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_114 VSS 1.22562f
C193 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_113 VSS 1.22562f
C194 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_112 VSS 1.22696f
C195 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_111 VSS 1.22562f
C196 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_110 VSS 1.22562f
C197 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_109 VSS 1.22562f
C198 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_108 VSS 1.22629f
C199 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_107 VSS 1.22696f
C200 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_106 VSS 1.22562f
C201 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_105 VSS 1.22562f
C202 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_104 VSS 1.22562f
C203 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_103 VSS 1.22629f
C204 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_102 VSS 1.22696f
C205 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_101 VSS 1.22562f
C206 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_100 VSS 1.22562f
C207 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 VSS 28.6559f
C208 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_98 VSS 1.22629f
C209 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_97 VSS 1.22562f
C210 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_96 VSS 1.22562f
C211 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_95 VSS 1.22562f
C212 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_94 VSS 1.22562f
C213 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_93 VSS 1.22629f
C214 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_92 VSS 1.22696f
C215 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_91 VSS 1.22562f
C216 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_90 VSS 1.22562f
C217 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_89 VSS 1.22629f
C218 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_88 VSS 1.22629f
C219 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_87 VSS 1.22562f
C220 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_86 VSS 1.22562f
C221 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_85 VSS 1.22562f
C222 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_84 VSS 1.22562f
C223 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_83 VSS 1.22629f
C224 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_82 VSS 1.22696f
C225 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_81 VSS 1.22562f
C226 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_80 VSS 1.22562f
C227 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_79 VSS 1.22562f
C228 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_78 VSS 1.22629f
C229 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_77 VSS 1.22562f
C230 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_76 VSS 1.22562f
C231 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_75 VSS 1.22562f
C232 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_74 VSS 1.22562f
C233 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_73 VSS 1.22629f
C234 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_72 VSS 1.22562f
C235 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_71 VSS 1.22562f
C236 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_70 VSS 1.22562f
C237 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_69 VSS 1.22562f
C238 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_68 VSS 1.22629f
C239 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_67 VSS 1.22696f
C240 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_66 VSS 1.22562f
C241 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_65 VSS 1.22562f
C242 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_64 VSS 1.22562f
C243 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_63 VSS 1.22629f
C244 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_62 VSS 1.22696f
C245 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_61 VSS 1.22562f
C246 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_60 VSS 1.22562f
C247 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_59 VSS 1.22562f
C248 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_58 VSS 1.22562f
C249 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_57 VSS 1.22696f
C250 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_56 VSS 1.22562f
C251 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_55 VSS 1.22562f
C252 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_54 VSS 1.22562f
C253 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_53 VSS 1.22629f
C254 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_52 VSS 1.22696f
C255 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_51 VSS 1.22562f
C256 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_50 VSS 1.22562f
C257 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_49 VSS 1.22562f
C258 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_48 VSS 1.22629f
C259 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_47 VSS 1.22562f
C260 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_46 VSS 1.22562f
C261 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_45 VSS 1.22562f
C262 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_44 VSS 1.22562f
C263 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_43 VSS 1.22629f
C264 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_42 VSS 1.22696f
C265 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_41 VSS 1.22562f
C266 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_40 VSS 1.22562f
C267 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_39 VSS 1.22562f
C268 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_38 VSS 1.22629f
C269 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_37 VSS 1.22562f
C270 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_35 VSS 1.22562f
C271 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_34 VSS 1.22562f
C272 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_33 VSS 1.22629f
C273 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_32 VSS 1.22696f
C274 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_31 VSS 1.22562f
C275 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_30 VSS 1.22562f
C276 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_29 VSS 1.22562f
C277 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_28 VSS 1.22629f
C278 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_27 VSS 1.22562f
C279 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_26 VSS 1.22562f
C280 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_25 VSS 1.22562f
C281 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_24 VSS 1.22562f
C282 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_23 VSS 1.22629f
C283 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_22 VSS 1.22696f
C284 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_21 VSS 1.22562f
C285 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_20 VSS 1.22562f
C286 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_19 VSS 1.22562f
C287 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_18 VSS 1.22629f
C288 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_16 VSS 1.22562f
C289 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_15 VSS 1.22562f
C290 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_14 VSS 1.22562f
C291 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_13 VSS 1.22562f
C292 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_12 VSS 1.22696f
C293 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_11 VSS 1.22562f
C294 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_10 VSS 1.22562f
C295 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_9 VSS 1.22562f
C296 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_8 VSS 1.22629f
C297 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_7 VSS 1.22562f
C298 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_6 VSS 1.22562f
C299 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_5 VSS 1.22562f
C300 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_4 VSS 1.22562f
C301 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_3 VSS 1.22896f
C302 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_2 VSS 1.22562f
C303 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_1 VSS 1.22562f
C304 resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_0 VSS 1.22562f
.ends

