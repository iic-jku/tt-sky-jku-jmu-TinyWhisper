magic
tech sky130A
magscale 1 2
timestamp 1757014995
<< nwell >>
rect -941 -1119 941 1119
<< pmoslvt >>
rect -745 -900 -545 900
rect -487 -900 -287 900
rect -229 -900 -29 900
rect 29 -900 229 900
rect 287 -900 487 900
rect 545 -900 745 900
<< pdiff >>
rect -803 888 -745 900
rect -803 -888 -791 888
rect -757 -888 -745 888
rect -803 -900 -745 -888
rect -545 888 -487 900
rect -545 -888 -533 888
rect -499 -888 -487 888
rect -545 -900 -487 -888
rect -287 888 -229 900
rect -287 -888 -275 888
rect -241 -888 -229 888
rect -287 -900 -229 -888
rect -29 888 29 900
rect -29 -888 -17 888
rect 17 -888 29 888
rect -29 -900 29 -888
rect 229 888 287 900
rect 229 -888 241 888
rect 275 -888 287 888
rect 229 -900 287 -888
rect 487 888 545 900
rect 487 -888 499 888
rect 533 -888 545 888
rect 487 -900 545 -888
rect 745 888 803 900
rect 745 -888 757 888
rect 791 -888 803 888
rect 745 -900 803 -888
<< pdiffc >>
rect -791 -888 -757 888
rect -533 -888 -499 888
rect -275 -888 -241 888
rect -17 -888 17 888
rect 241 -888 275 888
rect 499 -888 533 888
rect 757 -888 791 888
<< nsubdiff >>
rect -905 1049 -809 1083
rect 809 1049 905 1083
rect -905 987 -871 1049
rect 871 987 905 1049
rect -905 -1049 -871 -987
rect 871 -1049 905 -987
rect -905 -1083 -809 -1049
rect 809 -1083 905 -1049
<< nsubdiffcont >>
rect -809 1049 809 1083
rect -905 -987 -871 987
rect 871 -987 905 987
rect -809 -1083 809 -1049
<< poly >>
rect -745 981 -545 997
rect -745 947 -729 981
rect -561 947 -545 981
rect -745 900 -545 947
rect 545 981 745 997
rect 545 947 561 981
rect 729 947 745 981
rect -487 900 -287 945
rect -229 900 -29 945
rect 29 900 229 945
rect 287 900 487 945
rect 545 900 745 947
rect -745 -945 -545 -900
rect -487 -947 -287 -900
rect -487 -981 -471 -947
rect -303 -981 -287 -947
rect -487 -997 -287 -981
rect -229 -947 -29 -900
rect -229 -981 -213 -947
rect -45 -981 -29 -947
rect -229 -997 -29 -981
rect 29 -947 229 -900
rect 29 -981 45 -947
rect 213 -981 229 -947
rect 29 -997 229 -981
rect 287 -947 487 -900
rect 545 -945 745 -900
rect 287 -981 303 -947
rect 471 -981 487 -947
rect 287 -997 487 -981
<< polycont >>
rect -729 947 -561 981
rect 561 947 729 981
rect -471 -981 -303 -947
rect -213 -981 -45 -947
rect 45 -981 213 -947
rect 303 -981 471 -947
<< locali >>
rect -905 1049 -809 1083
rect 809 1049 905 1083
rect -905 987 -871 1049
rect 871 987 905 1049
rect -745 947 -729 981
rect -561 947 -545 981
rect 545 947 561 981
rect 729 947 745 981
rect -791 888 -757 904
rect -791 -904 -757 -888
rect -533 888 -499 904
rect -533 -904 -499 -888
rect -275 888 -241 904
rect -275 -904 -241 -888
rect -17 888 17 904
rect -17 -904 17 -888
rect 241 888 275 904
rect 241 -904 275 -888
rect 499 888 533 904
rect 499 -904 533 -888
rect 757 888 791 904
rect 757 -904 791 -888
rect -487 -981 -471 -947
rect -303 -981 -287 -947
rect -229 -981 -213 -947
rect -45 -981 -29 -947
rect 29 -981 45 -947
rect 213 -981 229 -947
rect 287 -981 303 -947
rect 471 -981 487 -947
rect -905 -1049 -871 -987
rect 871 -1049 905 -987
rect -905 -1083 -809 -1049
rect 809 -1083 905 -1049
<< viali >>
rect -729 947 -561 981
rect 561 947 729 981
rect -791 -888 -757 888
rect -533 -888 -499 888
rect -275 -888 -241 888
rect -17 -888 17 888
rect 241 -888 275 888
rect 499 -888 533 888
rect 757 -888 791 888
rect -471 -981 -303 -947
rect -213 -981 -45 -947
rect 45 -981 213 -947
rect 303 -981 471 -947
<< metal1 >>
rect -741 981 -549 987
rect -741 947 -729 981
rect -561 947 -549 981
rect -741 941 -549 947
rect 549 981 741 987
rect 549 947 561 981
rect 729 947 741 981
rect 549 941 741 947
rect -797 888 -751 900
rect -797 -888 -791 888
rect -757 -888 -751 888
rect -797 -900 -751 -888
rect -539 888 -493 900
rect -539 -888 -533 888
rect -499 -888 -493 888
rect -539 -900 -493 -888
rect -281 888 -235 900
rect -281 -888 -275 888
rect -241 -888 -235 888
rect -281 -900 -235 -888
rect -23 888 23 900
rect -23 -888 -17 888
rect 17 -888 23 888
rect -23 -900 23 -888
rect 235 888 281 900
rect 235 -888 241 888
rect 275 -888 281 888
rect 235 -900 281 -888
rect 493 888 539 900
rect 493 -888 499 888
rect 533 -888 539 888
rect 493 -900 539 -888
rect 751 888 797 900
rect 751 -888 757 888
rect 791 -888 797 888
rect 751 -900 797 -888
rect -483 -947 -291 -941
rect -483 -981 -471 -947
rect -303 -981 -291 -947
rect -483 -987 -291 -981
rect -225 -947 -33 -941
rect -225 -981 -213 -947
rect -45 -981 -33 -947
rect -225 -987 -33 -981
rect 33 -947 225 -941
rect 33 -981 45 -947
rect 213 -981 225 -947
rect 33 -987 225 -981
rect 291 -947 483 -941
rect 291 -981 303 -947
rect 471 -981 483 -947
rect 291 -987 483 -981
<< labels >>
rlabel nsubdiffcont 0 -1066 0 -1066 0 B
port 1 nsew
rlabel pdiffc -774 0 -774 0 0 D0
port 2 nsew
rlabel polycont -645 964 -645 964 0 G0
port 3 nsew
rlabel pdiffc -516 0 -516 0 0 S1
port 4 nsew
rlabel pdiffc -258 0 -258 0 0 D2
port 6 nsew
rlabel pdiffc 0 0 0 0 0 S3
port 8 nsew
rlabel pdiffc 258 0 258 0 0 D4
port 10 nsew
rlabel pdiffc 516 0 516 0 0 S5
port 12 nsew
rlabel polycont 645 964 645 964 0 G5
port 13 nsew
<< properties >>
string FIXED_BBOX -888 -1066 888 1066
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 9 l 1 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
