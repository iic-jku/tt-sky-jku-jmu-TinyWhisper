magic
tech sky130A
magscale 1 2
timestamp 1762641840
<< pwell >>
rect -1463 -310 1463 310
<< nmos >>
rect -1263 -100 -1233 100
rect -1167 -100 -1137 100
rect -1071 -100 -1041 100
rect -975 -100 -945 100
rect -879 -100 -849 100
rect -783 -100 -753 100
rect -687 -100 -657 100
rect -591 -100 -561 100
rect -495 -100 -465 100
rect -399 -100 -369 100
rect -303 -100 -273 100
rect -207 -100 -177 100
rect -111 -100 -81 100
rect -15 -100 15 100
rect 81 -100 111 100
rect 177 -100 207 100
rect 273 -100 303 100
rect 369 -100 399 100
rect 465 -100 495 100
rect 561 -100 591 100
rect 657 -100 687 100
rect 753 -100 783 100
rect 849 -100 879 100
rect 945 -100 975 100
rect 1041 -100 1071 100
rect 1137 -100 1167 100
rect 1233 -100 1263 100
<< ndiff >>
rect -1325 88 -1263 100
rect -1325 -88 -1313 88
rect -1279 -88 -1263 88
rect -1325 -100 -1263 -88
rect -1233 88 -1167 100
rect -1233 -88 -1217 88
rect -1183 -88 -1167 88
rect -1233 -100 -1167 -88
rect -1137 88 -1071 100
rect -1137 -88 -1121 88
rect -1087 -88 -1071 88
rect -1137 -100 -1071 -88
rect -1041 88 -975 100
rect -1041 -88 -1025 88
rect -991 -88 -975 88
rect -1041 -100 -975 -88
rect -945 88 -879 100
rect -945 -88 -929 88
rect -895 -88 -879 88
rect -945 -100 -879 -88
rect -849 88 -783 100
rect -849 -88 -833 88
rect -799 -88 -783 88
rect -849 -100 -783 -88
rect -753 88 -687 100
rect -753 -88 -737 88
rect -703 -88 -687 88
rect -753 -100 -687 -88
rect -657 88 -591 100
rect -657 -88 -641 88
rect -607 -88 -591 88
rect -657 -100 -591 -88
rect -561 88 -495 100
rect -561 -88 -545 88
rect -511 -88 -495 88
rect -561 -100 -495 -88
rect -465 88 -399 100
rect -465 -88 -449 88
rect -415 -88 -399 88
rect -465 -100 -399 -88
rect -369 88 -303 100
rect -369 -88 -353 88
rect -319 -88 -303 88
rect -369 -100 -303 -88
rect -273 88 -207 100
rect -273 -88 -257 88
rect -223 -88 -207 88
rect -273 -100 -207 -88
rect -177 88 -111 100
rect -177 -88 -161 88
rect -127 -88 -111 88
rect -177 -100 -111 -88
rect -81 88 -15 100
rect -81 -88 -65 88
rect -31 -88 -15 88
rect -81 -100 -15 -88
rect 15 88 81 100
rect 15 -88 31 88
rect 65 -88 81 88
rect 15 -100 81 -88
rect 111 88 177 100
rect 111 -88 127 88
rect 161 -88 177 88
rect 111 -100 177 -88
rect 207 88 273 100
rect 207 -88 223 88
rect 257 -88 273 88
rect 207 -100 273 -88
rect 303 88 369 100
rect 303 -88 319 88
rect 353 -88 369 88
rect 303 -100 369 -88
rect 399 88 465 100
rect 399 -88 415 88
rect 449 -88 465 88
rect 399 -100 465 -88
rect 495 88 561 100
rect 495 -88 511 88
rect 545 -88 561 88
rect 495 -100 561 -88
rect 591 88 657 100
rect 591 -88 607 88
rect 641 -88 657 88
rect 591 -100 657 -88
rect 687 88 753 100
rect 687 -88 703 88
rect 737 -88 753 88
rect 687 -100 753 -88
rect 783 88 849 100
rect 783 -88 799 88
rect 833 -88 849 88
rect 783 -100 849 -88
rect 879 88 945 100
rect 879 -88 895 88
rect 929 -88 945 88
rect 879 -100 945 -88
rect 975 88 1041 100
rect 975 -88 991 88
rect 1025 -88 1041 88
rect 975 -100 1041 -88
rect 1071 88 1137 100
rect 1071 -88 1087 88
rect 1121 -88 1137 88
rect 1071 -100 1137 -88
rect 1167 88 1233 100
rect 1167 -88 1183 88
rect 1217 -88 1233 88
rect 1167 -100 1233 -88
rect 1263 88 1325 100
rect 1263 -88 1279 88
rect 1313 -88 1325 88
rect 1263 -100 1325 -88
<< ndiffc >>
rect -1313 -88 -1279 88
rect -1217 -88 -1183 88
rect -1121 -88 -1087 88
rect -1025 -88 -991 88
rect -929 -88 -895 88
rect -833 -88 -799 88
rect -737 -88 -703 88
rect -641 -88 -607 88
rect -545 -88 -511 88
rect -449 -88 -415 88
rect -353 -88 -319 88
rect -257 -88 -223 88
rect -161 -88 -127 88
rect -65 -88 -31 88
rect 31 -88 65 88
rect 127 -88 161 88
rect 223 -88 257 88
rect 319 -88 353 88
rect 415 -88 449 88
rect 511 -88 545 88
rect 607 -88 641 88
rect 703 -88 737 88
rect 799 -88 833 88
rect 895 -88 929 88
rect 991 -88 1025 88
rect 1087 -88 1121 88
rect 1183 -88 1217 88
rect 1279 -88 1313 88
<< psubdiff >>
rect -1427 240 -1331 274
rect 1331 240 1427 274
rect -1427 178 -1393 240
rect 1393 178 1427 240
rect -1427 -240 -1393 -178
rect 1393 -240 1427 -178
rect -1427 -274 -1331 -240
rect 1331 -274 1427 -240
<< psubdiffcont >>
rect -1331 240 1331 274
rect -1427 -178 -1393 178
rect 1393 -178 1427 178
rect -1331 -274 1331 -240
<< poly >>
rect -1285 190 -925 225
rect -1285 155 -1260 190
rect -950 155 -925 190
rect -1285 120 -925 155
rect 925 190 1285 225
rect 925 155 950 190
rect 1260 155 1285 190
rect -1263 100 -1233 120
rect -1167 100 -1137 120
rect -1071 100 -1041 120
rect -975 100 -945 120
rect -879 100 -849 126
rect -783 100 -753 126
rect -687 100 -657 126
rect -591 100 -561 126
rect -495 100 -465 126
rect -399 100 -369 126
rect -303 100 -273 126
rect -207 100 -177 126
rect -111 100 -81 126
rect -15 100 15 126
rect 81 100 111 126
rect 177 100 207 126
rect 273 100 303 126
rect 369 100 399 126
rect 465 100 495 126
rect 561 100 591 126
rect 657 100 687 126
rect 753 100 783 126
rect 849 100 879 126
rect 925 120 1285 155
rect 945 100 975 120
rect 1041 100 1071 120
rect 1137 100 1167 120
rect 1233 100 1263 120
rect -1263 -126 -1233 -100
rect -1167 -126 -1137 -100
rect -1071 -126 -1041 -100
rect -975 -126 -945 -100
rect -879 -120 -849 -100
rect -783 -120 -753 -100
rect -687 -120 -657 -100
rect -591 -120 -561 -100
rect -495 -120 -465 -100
rect -399 -120 -369 -100
rect -303 -120 -273 -100
rect -207 -120 -177 -100
rect -111 -120 -81 -100
rect -15 -120 15 -100
rect 81 -120 111 -100
rect 177 -120 207 -100
rect 273 -120 303 -100
rect 369 -120 399 -100
rect 465 -120 495 -100
rect 561 -120 591 -100
rect 657 -120 687 -100
rect 753 -120 783 -100
rect 849 -120 879 -100
rect -900 -155 900 -120
rect 945 -126 975 -100
rect 1041 -126 1071 -100
rect 1137 -126 1167 -100
rect 1233 -126 1263 -100
rect -900 -190 -875 -155
rect 875 -190 900 -155
rect -900 -225 900 -190
<< polycont >>
rect -1260 155 -950 190
rect 950 155 1260 190
rect -875 -190 875 -155
<< locali >>
rect -1427 240 -1331 274
rect 1331 240 1427 274
rect -1427 178 -1393 240
rect -1280 190 -930 205
rect -1280 155 -1260 190
rect -950 155 -930 190
rect -1280 140 -930 155
rect 930 190 1280 205
rect 930 155 950 190
rect 1260 155 1280 190
rect 930 140 1280 155
rect 1393 178 1427 240
rect -1313 88 -1279 104
rect -1313 -104 -1279 -88
rect -1217 88 -1183 104
rect -1217 -104 -1183 -88
rect -1121 88 -1087 104
rect -1121 -104 -1087 -88
rect -1025 88 -991 104
rect -1025 -104 -991 -88
rect -929 88 -895 104
rect -929 -104 -895 -88
rect -833 88 -799 104
rect -833 -104 -799 -88
rect -737 88 -703 104
rect -737 -104 -703 -88
rect -641 88 -607 104
rect -641 -104 -607 -88
rect -545 88 -511 104
rect -545 -104 -511 -88
rect -449 88 -415 104
rect -449 -104 -415 -88
rect -353 88 -319 104
rect -353 -104 -319 -88
rect -257 88 -223 104
rect -257 -104 -223 -88
rect -161 88 -127 104
rect -161 -104 -127 -88
rect -65 88 -31 104
rect -65 -104 -31 -88
rect 31 88 65 104
rect 31 -104 65 -88
rect 127 88 161 104
rect 127 -104 161 -88
rect 223 88 257 104
rect 223 -104 257 -88
rect 319 88 353 104
rect 319 -104 353 -88
rect 415 88 449 104
rect 415 -104 449 -88
rect 511 88 545 104
rect 511 -104 545 -88
rect 607 88 641 104
rect 607 -104 641 -88
rect 703 88 737 104
rect 703 -104 737 -88
rect 799 88 833 104
rect 799 -104 833 -88
rect 895 88 929 104
rect 895 -104 929 -88
rect 991 88 1025 104
rect 991 -104 1025 -88
rect 1087 88 1121 104
rect 1087 -104 1121 -88
rect 1183 88 1217 104
rect 1183 -104 1217 -88
rect 1279 88 1313 104
rect 1279 -104 1313 -88
rect -1427 -240 -1393 -178
rect -895 -155 895 -140
rect -895 -190 -875 -155
rect 875 -190 895 -155
rect -895 -205 895 -190
rect 1393 -240 1427 -178
rect -1427 -274 -1331 -240
rect 1331 -274 1427 -240
<< viali >>
rect -1260 155 -950 190
rect 950 155 1260 190
rect -1313 -88 -1279 88
rect -1217 -88 -1183 88
rect -1121 -88 -1087 88
rect -1025 -88 -991 88
rect -929 -88 -895 88
rect -833 -88 -799 88
rect -737 -88 -703 88
rect -641 -88 -607 88
rect -545 -88 -511 88
rect -449 -88 -415 88
rect -353 -88 -319 88
rect -257 -88 -223 88
rect -161 -88 -127 88
rect -65 -88 -31 88
rect 31 -88 65 88
rect 127 -88 161 88
rect 223 -88 257 88
rect 319 -88 353 88
rect 415 -88 449 88
rect 511 -88 545 88
rect 607 -88 641 88
rect 703 -88 737 88
rect 799 -88 833 88
rect 895 -88 929 88
rect 991 -88 1025 88
rect 1087 -88 1121 88
rect 1183 -88 1217 88
rect 1279 -88 1313 88
rect -875 -190 875 -155
<< metal1 >>
rect -1280 190 -930 205
rect -1280 155 -1260 190
rect -950 155 -930 190
rect -1280 140 -930 155
rect 930 190 1280 205
rect 930 155 950 190
rect 1260 155 1280 190
rect 930 140 1280 155
rect -1319 88 -1273 100
rect -1319 -88 -1313 88
rect -1279 -88 -1273 88
rect -1319 -100 -1273 -88
rect -1223 88 -1177 100
rect -1223 -88 -1217 88
rect -1183 -88 -1177 88
rect -1223 -100 -1177 -88
rect -1127 88 -1081 100
rect -1127 -88 -1121 88
rect -1087 -88 -1081 88
rect -1127 -100 -1081 -88
rect -1031 88 -985 100
rect -1031 -88 -1025 88
rect -991 -88 -985 88
rect -1031 -100 -985 -88
rect -935 88 -889 100
rect -935 -88 -929 88
rect -895 -88 -889 88
rect -935 -100 -889 -88
rect -839 88 -793 100
rect -839 -88 -833 88
rect -799 -88 -793 88
rect -839 -100 -793 -88
rect -743 88 -697 100
rect -743 -88 -737 88
rect -703 -88 -697 88
rect -743 -100 -697 -88
rect -647 88 -601 100
rect -647 -88 -641 88
rect -607 -88 -601 88
rect -647 -100 -601 -88
rect -551 88 -505 100
rect -551 -88 -545 88
rect -511 -88 -505 88
rect -551 -100 -505 -88
rect -455 88 -409 100
rect -455 -88 -449 88
rect -415 -88 -409 88
rect -455 -100 -409 -88
rect -359 88 -313 100
rect -359 -88 -353 88
rect -319 -88 -313 88
rect -359 -100 -313 -88
rect -263 88 -217 100
rect -263 -88 -257 88
rect -223 -88 -217 88
rect -263 -100 -217 -88
rect -167 88 -121 100
rect -167 -88 -161 88
rect -127 -88 -121 88
rect -167 -100 -121 -88
rect -71 88 -25 100
rect -71 -88 -65 88
rect -31 -88 -25 88
rect -71 -100 -25 -88
rect 25 88 71 100
rect 25 -88 31 88
rect 65 -88 71 88
rect 25 -100 71 -88
rect 121 88 167 100
rect 121 -88 127 88
rect 161 -88 167 88
rect 121 -100 167 -88
rect 217 88 263 100
rect 217 -88 223 88
rect 257 -88 263 88
rect 217 -100 263 -88
rect 313 88 359 100
rect 313 -88 319 88
rect 353 -88 359 88
rect 313 -100 359 -88
rect 409 88 455 100
rect 409 -88 415 88
rect 449 -88 455 88
rect 409 -100 455 -88
rect 505 88 551 100
rect 505 -88 511 88
rect 545 -88 551 88
rect 505 -100 551 -88
rect 601 88 647 100
rect 601 -88 607 88
rect 641 -88 647 88
rect 601 -100 647 -88
rect 697 88 743 100
rect 697 -88 703 88
rect 737 -88 743 88
rect 697 -100 743 -88
rect 793 88 839 100
rect 793 -88 799 88
rect 833 -88 839 88
rect 793 -100 839 -88
rect 889 88 935 100
rect 889 -88 895 88
rect 929 -88 935 88
rect 889 -100 935 -88
rect 985 88 1031 100
rect 985 -88 991 88
rect 1025 -88 1031 88
rect 985 -100 1031 -88
rect 1081 88 1127 100
rect 1081 -88 1087 88
rect 1121 -88 1127 88
rect 1081 -100 1127 -88
rect 1177 88 1223 100
rect 1177 -88 1183 88
rect 1217 -88 1223 88
rect 1177 -100 1223 -88
rect 1273 88 1319 100
rect 1273 -88 1279 88
rect 1313 -88 1319 88
rect 1273 -100 1319 -88
rect -895 -155 895 -140
rect -895 -190 -875 -155
rect 875 -190 895 -155
rect -895 -205 895 -190
<< labels >>
rlabel psubdiffcont 0 -257 0 -257 0 B
port 1 nsew
rlabel ndiffc -1296 0 -1296 0 0 D0
port 2 nsew
rlabel ndiffc -1200 0 -1200 0 0 S1
port 4 nsew
rlabel ndiffc -1104 0 -1104 0 0 D2
port 6 nsew
rlabel ndiffc -1008 0 -1008 0 0 S3
port 8 nsew
rlabel ndiffc -912 0 -912 0 0 D4
port 10 nsew
rlabel poly -864 -155 -864 -155 0 G4
port 11 nsew
rlabel ndiffc -816 0 -816 0 0 S5
port 12 nsew
rlabel ndiffc -720 0 -720 0 0 D6
port 14 nsew
rlabel poly -672 -155 -672 -155 0 G6
port 15 nsew
rlabel ndiffc -624 0 -624 0 0 S7
port 16 nsew
rlabel ndiffc -528 0 -528 0 0 D8
port 18 nsew
rlabel poly -480 -155 -480 -155 0 G8
port 19 nsew
rlabel ndiffc -432 0 -432 0 0 S9
port 20 nsew
rlabel ndiffc -336 0 -336 0 0 D10
port 22 nsew
rlabel poly -288 -155 -288 -155 0 G10
port 23 nsew
rlabel ndiffc -240 0 -240 0 0 S11
port 24 nsew
rlabel ndiffc -144 0 -144 0 0 D12
port 26 nsew
rlabel poly -96 -155 -96 -155 0 G12
port 27 nsew
rlabel ndiffc -48 0 -48 0 0 S13
port 28 nsew
rlabel ndiffc 48 0 48 0 0 D14
port 30 nsew
rlabel poly 96 -155 96 -155 0 G14
port 31 nsew
rlabel ndiffc 144 0 144 0 0 S15
port 32 nsew
rlabel ndiffc 240 0 240 0 0 D16
port 34 nsew
rlabel poly 288 -155 288 -155 0 G16
port 35 nsew
rlabel ndiffc 336 0 336 0 0 S17
port 36 nsew
rlabel ndiffc 432 0 432 0 0 D18
port 38 nsew
rlabel poly 480 -155 480 -155 0 G18
port 39 nsew
rlabel ndiffc 528 0 528 0 0 S19
port 40 nsew
rlabel ndiffc 624 0 624 0 0 D20
port 42 nsew
rlabel poly 672 -155 672 -155 0 G20
port 43 nsew
rlabel ndiffc 720 0 720 0 0 S21
port 44 nsew
rlabel ndiffc 816 0 816 0 0 D22
port 46 nsew
rlabel poly 864 -155 864 -155 0 G22
port 47 nsew
rlabel ndiffc 912 0 912 0 0 S23
port 48 nsew
rlabel poly 960 155 960 155 0 G23
port 49 nsew
rlabel ndiffc 1008 0 1008 0 0 D24
port 50 nsew
rlabel ndiffc 1104 0 1104 0 0 S25
port 52 nsew
rlabel poly 1152 155 1152 155 0 G25
port 53 nsew
rlabel ndiffc 1200 0 1200 0 0 D26
port 54 nsew
rlabel ndiffc 1296 0 1296 0 0 S26
port 55 nsew
rlabel poly -960 155 -960 155 0 G3
port 9 nsew
rlabel poly -1152 155 -1152 155 0 G1
port 5 nsew
<< properties >>
string FIXED_BBOX -1410 -257 1410 257
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.15 m 1 nf 27 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
