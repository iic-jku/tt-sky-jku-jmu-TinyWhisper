magic
tech sky130A
magscale 1 2
timestamp 1762093820
<< metal1 >>
rect 4848 9580 5253 9586
rect 4214 9175 4220 9580
rect 4625 9175 4631 9580
rect 4848 9175 6246 9580
rect 4848 9169 5253 9175
rect 4234 6184 4240 6294
rect 4350 6184 4356 6294
rect 6564 2243 6969 4535
rect 6564 1838 19047 2243
rect 18642 1735 19047 1838
rect 18641 1729 19048 1735
rect 18641 1316 19048 1322
<< via1 >>
rect 4220 9175 4625 9580
rect 4240 6184 4350 6294
rect 18641 1322 19048 1729
<< metal2 >>
rect 4220 9580 4625 9586
rect 2403 9175 4220 9580
rect 2403 8493 2808 9175
rect 4220 9169 4625 9175
rect 2403 8089 2808 8098
rect 4240 6294 4350 6300
rect 3310 6184 4240 6294
rect 3311 1304 3419 6184
rect 4240 6178 4350 6184
rect 18635 1322 18641 1729
rect 19048 1322 19054 1729
rect 18641 1313 19048 1322
rect 3311 1196 12551 1304
rect 12649 1196 12658 1304
<< via2 >>
rect 2403 8098 2808 8493
rect 18641 1322 19048 1719
rect 12551 1196 12649 1304
<< metal3 >>
rect 33607 8645 33613 9580
rect 34546 8645 34552 9580
rect 2398 8496 2813 8502
rect 2398 8087 2813 8093
rect 2398 5569 2404 5972
rect 2807 5569 2813 5972
rect 7585 2380 8506 7111
rect 32825 3165 33745 5050
rect 26115 2245 33745 3165
rect 26115 2098 27035 2245
rect 18636 1722 19053 1728
rect 18636 1311 19053 1317
rect 12546 1304 12654 1309
rect 14946 1304 15054 1308
rect 12546 1196 12551 1304
rect 12649 1302 15054 1304
rect 12649 1196 14946 1302
rect 12546 1191 12654 1196
rect 14946 1190 15054 1196
rect 26115 1174 27035 1180
<< via3 >>
rect 33613 8645 34546 9580
rect 2398 8493 2813 8496
rect 2398 8098 2403 8493
rect 2403 8098 2808 8493
rect 2808 8098 2813 8493
rect 2398 8093 2813 8098
rect 2404 5569 2807 5972
rect 18636 1719 19053 1722
rect 18636 1322 18641 1719
rect 18641 1322 19048 1719
rect 19048 1322 19053 1719
rect 18636 1317 19053 1322
rect 14946 1196 15054 1302
rect 26115 1180 27035 2098
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 44952 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 200 1000 600 44152
rect 800 1000 1200 44152
rect 33612 9580 34547 9581
rect 33612 8645 33613 9580
rect 34546 8645 34547 9580
rect 2397 8496 2814 8497
rect 2397 8093 2398 8496
rect 2813 8093 2814 8496
rect 2397 8092 2814 8093
rect 2403 5972 2808 8092
rect 2403 5945 2404 5972
rect 2398 5569 2404 5945
rect 2807 5569 2808 5972
rect 2398 5568 2808 5569
rect 2398 2707 2803 5568
rect 2398 2303 22922 2707
rect 18639 1723 19049 1724
rect 18635 1722 19054 1723
rect 18635 1317 18636 1722
rect 19053 1317 19054 1722
rect 18635 1316 19054 1317
rect 14945 1302 15055 1303
rect 14945 1196 14946 1302
rect 15054 1196 15055 1302
rect 14945 1195 15055 1196
rect 14946 200 15054 1195
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18639 25 19049 1316
rect 22518 58 22922 2303
rect 33612 2148 34547 8645
rect 26114 2098 27036 2099
rect 26114 1180 26115 2098
rect 27035 1180 27036 2098
rect 26114 1179 27036 1180
rect 29953 1213 34547 2148
rect 18770 0 18950 25
rect 22634 0 22814 58
rect 26115 55 27035 1179
rect 29953 78 30888 1213
rect 26498 0 26678 55
rect 30362 0 30542 78
use third_order_mfb_lp_filter  third_order_mfb_lp_filter_0 /foss/designs/tt-sky-jku-jmu-TinyWhisper/mag/third_order_mfb_lp_filter
timestamp 1762090404
transform 1 0 6325 0 1 3030
box -2685 40 28500 7610
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 66976 45152
<< end >>
