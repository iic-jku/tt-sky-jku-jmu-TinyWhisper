magic
tech sky130A
magscale 1 2
timestamp 1761785752
<< locali >>
rect -30 8175 75 8190
rect -30 8080 -15 8175
rect 60 8080 75 8175
rect -30 8065 75 8080
rect -30 2335 75 2350
rect -30 2240 -15 2335
rect 60 2240 75 2335
rect -30 2225 75 2240
<< viali >>
rect -15 8080 60 8175
rect -15 2240 60 2335
<< metal1 >>
rect 6120 8985 16830 8995
rect 6120 8925 16720 8985
rect 16820 8925 16830 8985
rect 6120 8915 16830 8925
rect 6120 8330 6345 8915
rect 16745 8330 16830 8735
rect -65 8175 75 8190
rect -65 8080 -15 8175
rect 60 8080 75 8175
rect -65 8065 75 8080
rect -65 7530 200 7935
rect 2965 7315 3190 7935
rect 16545 7315 16665 7935
rect 16710 7500 16830 7935
rect 23115 7530 23150 7935
rect 16710 7435 16725 7500
rect 16815 7435 16830 7500
rect 16710 7420 16830 7435
rect -65 2485 200 2890
rect 2970 2485 3185 3105
rect 16545 2485 16665 3105
rect 16710 2985 16830 3000
rect 16710 2920 16725 2985
rect 16815 2920 16830 2985
rect 16710 2485 16830 2920
rect 23115 2485 23150 2890
rect -65 2335 75 2350
rect -65 2240 -15 2335
rect 60 2240 75 2335
rect -65 2225 75 2240
rect 6120 1505 6340 2090
rect 16745 1685 16830 2090
rect 6120 1495 16830 1505
rect 6120 1435 16720 1495
rect 16820 1435 16830 1495
rect 6120 1425 16830 1435
<< via1 >>
rect 16720 8925 16820 8985
rect 16725 7435 16815 7500
rect 16725 2920 16815 2985
rect 16720 1435 16820 1495
<< metal2 >>
rect 16710 8985 16830 8995
rect 16710 8925 16720 8985
rect 16820 8925 16830 8985
rect 16710 7500 16830 8925
rect 16710 7435 16725 7500
rect 16815 7435 16830 7500
rect 16710 7420 16830 7435
rect 16710 2985 16830 3000
rect 16710 2920 16725 2985
rect 16815 2920 16830 2985
rect 16710 1495 16830 2920
rect 16710 1435 16720 1495
rect 16820 1435 16830 1495
rect 16710 1425 16830 1435
use resistors_n  resistors_n_0
timestamp 1757114530
transform 1 0 -165 0 1 -5845
box 100 7350 23315 8914
use resistors_p  resistors_p_0
timestamp 1757114131
transform 1 0 0 0 1 0
box -65 7350 23150 8914
<< end >>
