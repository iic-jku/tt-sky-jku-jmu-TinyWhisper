magic
tech sky130A
magscale 1 2
timestamp 1762641840
<< nwell >>
rect 15 670 4795 1710
rect 15 -1190 4795 -150
<< locali >>
rect 15 1865 4795 1880
rect 15 1755 30 1865
rect 4780 1755 4795 1865
rect 15 1640 4795 1755
rect 665 670 1005 1640
rect 1585 670 1925 1640
rect 2505 670 2845 1640
rect 3425 670 3765 1640
rect 665 70 1005 620
rect 1585 70 1925 620
rect 2505 70 2845 620
rect 3425 70 3765 620
rect 15 0 4795 70
rect 15 -220 4795 -150
rect 470 -1190 1005 -220
rect 1585 -1190 1925 -220
rect 2505 -1190 2845 -220
rect 3425 -1190 3765 -220
rect 470 -1790 1005 -1240
rect 1585 -1790 1925 -1240
rect 2505 -1790 2845 -1240
rect 3425 -1790 3765 -1240
rect 15 -1905 4795 -1790
rect 15 -2015 30 -1905
rect 4780 -2015 4795 -1905
rect 15 -2030 4795 -2015
<< viali >>
rect 30 1755 4780 1865
rect 30 -2015 4780 -1905
<< metal1 >>
rect 15 1865 4795 1880
rect 15 1755 30 1865
rect 4780 1755 4795 1865
rect 15 1640 4795 1755
rect 1600 1465 1910 1640
rect 1600 915 1700 1465
rect 1810 915 1910 1465
rect 1600 890 1910 915
rect 2520 1465 2830 1640
rect 2520 915 2620 1465
rect 2730 915 2830 1465
rect 2520 890 2830 915
rect -195 585 5 705
rect 785 695 920 705
rect 785 595 795 695
rect 875 595 920 695
rect 785 585 920 595
rect 1705 695 1855 705
rect 3545 695 3695 705
rect 1705 595 1715 695
rect 1795 595 1855 695
rect 3545 595 3555 695
rect 3635 595 3695 695
rect 1705 585 1855 595
rect 3545 585 3695 595
rect -195 -1155 -75 585
rect 680 385 990 410
rect 680 70 780 385
rect 15 25 780 70
rect 890 70 990 385
rect 3440 385 3750 410
rect 3440 70 3540 385
rect 890 25 3540 70
rect 3650 70 3750 385
rect 3650 25 4795 70
rect 15 0 4795 25
rect 15 -220 4795 -150
rect 1600 -395 1910 -220
rect 1600 -945 1700 -395
rect 1810 -945 1910 -395
rect 1600 -970 1910 -945
rect 2520 -395 2830 -220
rect 2520 -945 2620 -395
rect 2730 -945 2830 -395
rect 2520 -970 2830 -945
rect 470 -1030 545 -1020
rect 470 -1095 480 -1030
rect 535 -1095 545 -1030
rect -195 -1275 0 -1155
rect 470 -1450 545 -1095
rect 785 -1165 935 -1155
rect 785 -1265 795 -1165
rect 875 -1265 935 -1165
rect 785 -1275 935 -1265
rect 1705 -1165 1855 -1155
rect 3545 -1165 3695 -1155
rect 1705 -1265 1715 -1165
rect 1795 -1265 1855 -1165
rect 3545 -1265 3555 -1165
rect 3635 -1265 3695 -1165
rect 1705 -1275 1855 -1265
rect 3545 -1275 3695 -1265
rect 470 -1475 990 -1450
rect 470 -1790 780 -1475
rect 15 -1835 780 -1790
rect 890 -1790 990 -1475
rect 3440 -1475 3750 -1450
rect 3440 -1790 3540 -1475
rect 890 -1835 3540 -1790
rect 3650 -1790 3750 -1475
rect 3650 -1835 4795 -1790
rect 15 -1905 4795 -1835
rect 15 -2015 30 -1905
rect 4780 -2015 4795 -1905
rect 15 -2030 4795 -2015
<< via1 >>
rect 1700 915 1810 1465
rect 2620 915 2730 1465
rect 795 595 875 695
rect 1715 595 1795 695
rect 2050 595 2190 695
rect 2970 595 3110 695
rect 3555 595 3635 695
rect 780 25 890 385
rect 3540 25 3650 385
rect 205 -320 355 -265
rect 25 -960 80 -375
rect 1700 -945 1810 -395
rect 2620 -945 2730 -395
rect 480 -1095 535 -1030
rect 795 -1265 875 -1165
rect 1715 -1265 1795 -1165
rect 2050 -1265 2190 -1165
rect 2970 -1265 3110 -1165
rect 3555 -1265 3635 -1165
rect 780 -1835 890 -1475
rect 3540 -1835 3650 -1475
<< metal2 >>
rect 1690 1465 1820 1475
rect 1690 915 1700 1465
rect 1810 915 1820 1465
rect 1690 905 1820 915
rect 2610 1465 2740 1475
rect 2610 915 2620 1465
rect 2730 915 2740 1465
rect 2610 905 2740 915
rect 750 695 885 705
rect 750 595 795 695
rect 875 595 885 695
rect 750 585 885 595
rect 1655 695 1805 705
rect 1655 595 1715 695
rect 1795 595 1805 695
rect 1655 585 1805 595
rect 2040 695 2200 705
rect 2960 695 3120 705
rect 2040 595 2050 695
rect 2190 595 2200 695
rect 2960 595 2970 695
rect 3110 595 3120 695
rect 2040 585 2200 595
rect 2960 585 3120 595
rect 3510 695 3645 705
rect 3510 595 3555 695
rect 3635 595 3645 695
rect 3510 585 3645 595
rect 4795 585 5005 705
rect 770 385 900 395
rect 770 25 780 385
rect 890 25 900 385
rect 770 15 900 25
rect 3530 385 3660 395
rect 3530 25 3540 385
rect 3650 25 3660 385
rect 3530 15 3660 25
rect 2295 -20 3170 -10
rect 2295 -130 2305 -20
rect 2430 -130 3035 -20
rect 3160 -130 3170 -20
rect 2295 -140 3170 -130
rect 195 -265 545 -255
rect 195 -320 205 -265
rect 355 -320 545 -265
rect 195 -330 545 -320
rect 15 -375 90 -365
rect 15 -960 25 -375
rect 80 -960 90 -375
rect 15 -1685 90 -960
rect 470 -1030 545 -330
rect 1690 -395 1820 -385
rect 1690 -945 1700 -395
rect 1810 -945 1820 -395
rect 1690 -955 1820 -945
rect 2610 -395 2740 -385
rect 2610 -945 2620 -395
rect 2730 -945 2740 -395
rect 2610 -955 2740 -945
rect 470 -1095 480 -1030
rect 535 -1095 545 -1030
rect 470 -1105 545 -1095
rect 485 -1165 885 -1155
rect 485 -1265 795 -1165
rect 875 -1265 885 -1165
rect 485 -1275 885 -1265
rect 1670 -1165 1805 -1155
rect 1670 -1265 1715 -1165
rect 1795 -1265 1805 -1165
rect 1670 -1275 1805 -1265
rect 2040 -1165 2200 -1155
rect 2960 -1165 3120 -1155
rect 2040 -1265 2050 -1165
rect 2190 -1265 2200 -1165
rect 2960 -1265 2970 -1165
rect 3110 -1265 3120 -1165
rect 2040 -1275 2200 -1265
rect 2960 -1275 3120 -1265
rect 3510 -1165 3645 -1155
rect 3510 -1265 3555 -1165
rect 3635 -1265 3645 -1165
rect 3510 -1275 3645 -1265
rect 4795 -1275 5005 -1155
rect 770 -1475 900 -1465
rect 15 -1760 365 -1685
rect 770 -1835 780 -1475
rect 890 -1835 900 -1475
rect 770 -1845 900 -1835
rect 3530 -1475 3660 -1465
rect 3530 -1835 3540 -1475
rect 3650 -1835 3660 -1475
rect 3530 -1845 3660 -1835
<< via2 >>
rect 1700 915 1810 1465
rect 2620 915 2730 1465
rect 2050 595 2190 695
rect 2305 595 2430 695
rect 2970 595 3110 695
rect 780 25 890 385
rect 3540 25 3650 385
rect 2305 -130 2430 -20
rect 3035 -130 3160 -20
rect 1700 -945 1810 -395
rect 2620 -945 2730 -395
rect 2050 -1265 2190 -1165
rect 2305 -1265 2430 -1165
rect 2970 -1265 3110 -1165
rect 780 -1835 890 -1475
rect 3540 -1835 3650 -1475
<< metal3 >>
rect 1990 1565 3055 1710
rect 1600 1465 1910 1490
rect 1600 915 1700 1465
rect 1810 915 1910 1465
rect 680 385 990 410
rect 680 25 780 385
rect 890 25 990 385
rect 680 -1475 990 25
rect 1600 -395 1910 915
rect 1600 -945 1700 -395
rect 1810 -945 1910 -395
rect 1600 -970 1910 -945
rect 1990 705 2135 1565
rect 2520 1465 2830 1490
rect 2520 915 2620 1465
rect 2730 915 2830 1465
rect 1990 695 2200 705
rect 1990 595 2050 695
rect 2190 595 2200 695
rect 1990 585 2200 595
rect 2295 695 2440 705
rect 2295 595 2305 695
rect 2430 595 2440 695
rect 1990 -915 2135 585
rect 2295 -20 2440 595
rect 2295 -130 2305 -20
rect 2430 -130 2440 -20
rect 2295 -140 2440 -130
rect 2520 -395 2830 915
rect 2910 705 3055 1565
rect 2910 695 3120 705
rect 2910 595 2970 695
rect 3110 595 3120 695
rect 2910 585 3120 595
rect 3440 385 3750 410
rect 3440 25 3540 385
rect 3650 25 3750 385
rect 1990 -1060 2415 -915
rect 2520 -945 2620 -395
rect 2730 -945 2830 -395
rect 2520 -970 2830 -945
rect 3025 -20 3170 -10
rect 3025 -130 3035 -20
rect 3160 -130 3170 -20
rect 2295 -1155 2415 -1060
rect 3025 -1155 3170 -130
rect 680 -1835 780 -1475
rect 890 -1835 990 -1475
rect 1990 -1165 2200 -1155
rect 1990 -1265 2050 -1165
rect 2190 -1265 2200 -1165
rect 1990 -1275 2200 -1265
rect 2295 -1165 2440 -1155
rect 2295 -1265 2305 -1165
rect 2430 -1265 2440 -1165
rect 2295 -1275 2440 -1265
rect 2960 -1165 3170 -1155
rect 2960 -1265 2970 -1165
rect 3110 -1265 3170 -1165
rect 2960 -1275 3170 -1265
rect 1990 -1370 2135 -1275
rect 3025 -1370 3170 -1275
rect 1990 -1515 3170 -1370
rect 3440 -1475 3750 25
rect 680 -1860 990 -1835
rect 3440 -1835 3540 -1475
rect 3650 -1835 3750 -1475
rect 3440 -1860 3750 -1835
use inverter_NF1  inverter_NF1_0 inverter/inverter_NF1
timestamp 1762641840
transform 1 0 1910 0 1 725
box -70 -725 680 985
use inverter_NF1  inverter_NF1_1
timestamp 1762641840
transform 1 0 1910 0 1 -1135
box -70 -725 680 985
use inverter_NF2  inverter_NF2_0 inverter/inverter_NF2
timestamp 1762641840
transform 1 0 70 0 1 725
box -70 -725 680 985
use inverter_NF2  inverter_NF2_1
timestamp 1762641840
transform 1 0 990 0 1 725
box -70 -725 680 985
use inverter_NF2  inverter_NF2_2
timestamp 1762641840
transform 1 0 990 0 1 -1135
box -70 -725 680 985
use inverter_NF2  inverter_NF2_3
timestamp 1762641840
transform 1 0 2830 0 1 -1135
box -70 -725 680 985
use inverter_NF2  inverter_NF2_4
timestamp 1762641840
transform 1 0 2830 0 1 725
box -70 -725 680 985
use inverter_NF6  inverter_NF6_0 inverter/inverter_NF6
timestamp 1762641840
transform 1 0 3750 0 1 725
box -70 -725 1060 985
use inverter_NF6  inverter_NF6_1
timestamp 1762641840
transform 1 0 3750 0 1 -1135
box -70 -725 1060 985
use transmission_gate_wo_dummy  transmission_gate_wo_dummy_0 transmission_gate_wo_dummy
timestamp 1762641840
transform 1 0 70 0 1 -1135
box -70 -725 490 986
<< labels >>
flabel metal2 4905 645 4905 645 0 FreeSans 480 0 0 0 vout_LO
port 11 nsew
flabel metal2 4900 -1215 4900 -1215 0 FreeSans 480 0 0 0 vout_LO_inv
port 13 nsew
flabel space 3890 -1215 3890 -1215 0 FreeSans 320 0 0 0 inv_scale
flabel via2 2070 -1220 2070 -1220 0 FreeSans 320 0 0 0 inv_cross
flabel via2 2065 650 2065 650 0 FreeSans 320 0 0 0 buf_cross
flabel metal1 -135 -235 -135 -235 0 FreeSans 480 0 0 0 vin_LO
port 9 nsew
flabel viali 2210 1810 2210 1810 0 FreeSans 800 0 0 0 VDD
port 17 nsew
flabel space 3915 645 3915 645 0 FreeSans 320 0 0 0 buf_scale
flabel viali 2210 -1975 2210 -1975 0 FreeSans 800 0 0 0 VSS
port 15 nsew
<< end >>
