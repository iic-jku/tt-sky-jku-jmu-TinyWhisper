magic
tech sky130A
magscale 1 2
timestamp 1762641840
<< nwell >>
rect -1463 -519 1463 519
<< pmos >>
rect -1263 -300 -1233 300
rect -1167 -300 -1137 300
rect -1071 -300 -1041 300
rect -975 -300 -945 300
rect -879 -300 -849 300
rect -783 -300 -753 300
rect -687 -300 -657 300
rect -591 -300 -561 300
rect -495 -300 -465 300
rect -399 -300 -369 300
rect -303 -300 -273 300
rect -207 -300 -177 300
rect -111 -300 -81 300
rect -15 -300 15 300
rect 81 -300 111 300
rect 177 -300 207 300
rect 273 -300 303 300
rect 369 -300 399 300
rect 465 -300 495 300
rect 561 -300 591 300
rect 657 -300 687 300
rect 753 -300 783 300
rect 849 -300 879 300
rect 945 -300 975 300
rect 1041 -300 1071 300
rect 1137 -300 1167 300
rect 1233 -300 1263 300
<< pdiff >>
rect -1325 288 -1263 300
rect -1325 -288 -1313 288
rect -1279 -288 -1263 288
rect -1325 -300 -1263 -288
rect -1233 288 -1167 300
rect -1233 -288 -1217 288
rect -1183 -288 -1167 288
rect -1233 -300 -1167 -288
rect -1137 288 -1071 300
rect -1137 -288 -1121 288
rect -1087 -288 -1071 288
rect -1137 -300 -1071 -288
rect -1041 288 -975 300
rect -1041 -288 -1025 288
rect -991 -288 -975 288
rect -1041 -300 -975 -288
rect -945 288 -879 300
rect -945 -288 -929 288
rect -895 -288 -879 288
rect -945 -300 -879 -288
rect -849 288 -783 300
rect -849 -288 -833 288
rect -799 -288 -783 288
rect -849 -300 -783 -288
rect -753 288 -687 300
rect -753 -288 -737 288
rect -703 -288 -687 288
rect -753 -300 -687 -288
rect -657 288 -591 300
rect -657 -288 -641 288
rect -607 -288 -591 288
rect -657 -300 -591 -288
rect -561 288 -495 300
rect -561 -288 -545 288
rect -511 -288 -495 288
rect -561 -300 -495 -288
rect -465 288 -399 300
rect -465 -288 -449 288
rect -415 -288 -399 288
rect -465 -300 -399 -288
rect -369 288 -303 300
rect -369 -288 -353 288
rect -319 -288 -303 288
rect -369 -300 -303 -288
rect -273 288 -207 300
rect -273 -288 -257 288
rect -223 -288 -207 288
rect -273 -300 -207 -288
rect -177 288 -111 300
rect -177 -288 -161 288
rect -127 -288 -111 288
rect -177 -300 -111 -288
rect -81 288 -15 300
rect -81 -288 -65 288
rect -31 -288 -15 288
rect -81 -300 -15 -288
rect 15 288 81 300
rect 15 -288 31 288
rect 65 -288 81 288
rect 15 -300 81 -288
rect 111 288 177 300
rect 111 -288 127 288
rect 161 -288 177 288
rect 111 -300 177 -288
rect 207 288 273 300
rect 207 -288 223 288
rect 257 -288 273 288
rect 207 -300 273 -288
rect 303 288 369 300
rect 303 -288 319 288
rect 353 -288 369 288
rect 303 -300 369 -288
rect 399 288 465 300
rect 399 -288 415 288
rect 449 -288 465 288
rect 399 -300 465 -288
rect 495 288 561 300
rect 495 -288 511 288
rect 545 -288 561 288
rect 495 -300 561 -288
rect 591 288 657 300
rect 591 -288 607 288
rect 641 -288 657 288
rect 591 -300 657 -288
rect 687 288 753 300
rect 687 -288 703 288
rect 737 -288 753 288
rect 687 -300 753 -288
rect 783 288 849 300
rect 783 -288 799 288
rect 833 -288 849 288
rect 783 -300 849 -288
rect 879 288 945 300
rect 879 -288 895 288
rect 929 -288 945 288
rect 879 -300 945 -288
rect 975 288 1041 300
rect 975 -288 991 288
rect 1025 -288 1041 288
rect 975 -300 1041 -288
rect 1071 288 1137 300
rect 1071 -288 1087 288
rect 1121 -288 1137 288
rect 1071 -300 1137 -288
rect 1167 288 1233 300
rect 1167 -288 1183 288
rect 1217 -288 1233 288
rect 1167 -300 1233 -288
rect 1263 288 1325 300
rect 1263 -288 1279 288
rect 1313 -288 1325 288
rect 1263 -300 1325 -288
<< pdiffc >>
rect -1313 -288 -1279 288
rect -1217 -288 -1183 288
rect -1121 -288 -1087 288
rect -1025 -288 -991 288
rect -929 -288 -895 288
rect -833 -288 -799 288
rect -737 -288 -703 288
rect -641 -288 -607 288
rect -545 -288 -511 288
rect -449 -288 -415 288
rect -353 -288 -319 288
rect -257 -288 -223 288
rect -161 -288 -127 288
rect -65 -288 -31 288
rect 31 -288 65 288
rect 127 -288 161 288
rect 223 -288 257 288
rect 319 -288 353 288
rect 415 -288 449 288
rect 511 -288 545 288
rect 607 -288 641 288
rect 703 -288 737 288
rect 799 -288 833 288
rect 895 -288 929 288
rect 991 -288 1025 288
rect 1087 -288 1121 288
rect 1183 -288 1217 288
rect 1279 -288 1313 288
<< nsubdiff >>
rect -1427 449 -1331 483
rect 1331 449 1427 483
rect -1427 387 -1393 449
rect 1393 387 1427 449
rect -1427 -449 -1393 -387
rect 1393 -449 1427 -387
rect -1427 -483 -1331 -449
rect 1331 -483 1427 -449
<< nsubdiffcont >>
rect -1331 449 1331 483
rect -1427 -387 -1393 387
rect 1393 -387 1427 387
rect -1331 -483 1331 -449
<< poly >>
rect -1285 395 -925 430
rect -1285 360 -1260 395
rect -950 360 -925 395
rect -1285 325 -925 360
rect 925 395 1285 430
rect 925 360 950 395
rect 1260 360 1285 395
rect -1263 300 -1233 325
rect -1167 300 -1137 325
rect -1071 300 -1041 325
rect -975 300 -945 325
rect -879 300 -849 326
rect -783 300 -753 326
rect -687 300 -657 326
rect -591 300 -561 326
rect -495 300 -465 326
rect -399 300 -369 326
rect -303 300 -273 326
rect -207 300 -177 326
rect -111 300 -81 326
rect -15 300 15 326
rect 81 300 111 326
rect 177 300 207 326
rect 273 300 303 326
rect 369 300 399 326
rect 465 300 495 326
rect 561 300 591 326
rect 657 300 687 326
rect 753 300 783 326
rect 849 300 879 326
rect 925 325 1285 360
rect 945 300 975 325
rect 1041 300 1071 325
rect 1137 300 1167 325
rect 1233 300 1263 325
rect -1263 -326 -1233 -300
rect -1167 -326 -1137 -300
rect -1071 -326 -1041 -300
rect -975 -326 -945 -300
rect -879 -325 -849 -300
rect -783 -325 -753 -300
rect -687 -325 -657 -300
rect -591 -325 -561 -300
rect -495 -325 -465 -300
rect -399 -325 -369 -300
rect -303 -325 -273 -300
rect -207 -325 -177 -300
rect -111 -325 -81 -300
rect -15 -325 15 -300
rect 81 -325 111 -300
rect 177 -325 207 -300
rect 273 -325 303 -300
rect 369 -325 399 -300
rect 465 -325 495 -300
rect 561 -325 591 -300
rect 657 -325 687 -300
rect 753 -325 783 -300
rect 849 -325 879 -300
rect -900 -360 900 -325
rect 945 -326 975 -300
rect 1041 -326 1071 -300
rect 1137 -326 1167 -300
rect 1233 -326 1263 -300
rect -900 -395 -875 -360
rect 875 -395 900 -360
rect -900 -430 900 -395
<< polycont >>
rect -1260 360 -950 395
rect 950 360 1260 395
rect -875 -395 875 -360
<< locali >>
rect -1427 449 -1331 483
rect 1331 449 1427 483
rect -1427 387 -1393 449
rect -1280 395 -930 415
rect -1280 360 -1260 395
rect -950 360 -930 395
rect -1280 340 -930 360
rect 930 395 1280 415
rect 930 360 950 395
rect 1260 360 1280 395
rect 930 340 1280 360
rect 1393 387 1427 449
rect -1313 288 -1279 304
rect -1313 -304 -1279 -288
rect -1217 288 -1183 304
rect -1217 -304 -1183 -288
rect -1121 288 -1087 304
rect -1121 -304 -1087 -288
rect -1025 288 -991 304
rect -1025 -304 -991 -288
rect -929 288 -895 304
rect -929 -304 -895 -288
rect -833 288 -799 304
rect -833 -304 -799 -288
rect -737 288 -703 304
rect -737 -304 -703 -288
rect -641 288 -607 304
rect -641 -304 -607 -288
rect -545 288 -511 304
rect -545 -304 -511 -288
rect -449 288 -415 304
rect -449 -304 -415 -288
rect -353 288 -319 304
rect -353 -304 -319 -288
rect -257 288 -223 304
rect -257 -304 -223 -288
rect -161 288 -127 304
rect -161 -304 -127 -288
rect -65 288 -31 304
rect -65 -304 -31 -288
rect 31 288 65 304
rect 31 -304 65 -288
rect 127 288 161 304
rect 127 -304 161 -288
rect 223 288 257 304
rect 223 -304 257 -288
rect 319 288 353 304
rect 319 -304 353 -288
rect 415 288 449 304
rect 415 -304 449 -288
rect 511 288 545 304
rect 511 -304 545 -288
rect 607 288 641 304
rect 607 -304 641 -288
rect 703 288 737 304
rect 703 -304 737 -288
rect 799 288 833 304
rect 799 -304 833 -288
rect 895 288 929 304
rect 895 -304 929 -288
rect 991 288 1025 304
rect 991 -304 1025 -288
rect 1087 288 1121 304
rect 1087 -304 1121 -288
rect 1183 288 1217 304
rect 1183 -304 1217 -288
rect 1279 288 1313 304
rect 1279 -304 1313 -288
rect -1427 -449 -1393 -387
rect -895 -360 895 -340
rect -895 -395 -875 -360
rect 875 -395 895 -360
rect -895 -415 895 -395
rect 1393 -449 1427 -387
rect -1427 -483 -1331 -449
rect 1331 -483 1427 -449
<< viali >>
rect -1260 360 -950 395
rect 950 360 1260 395
rect -1313 -288 -1279 288
rect -1217 -288 -1183 288
rect -1121 -288 -1087 288
rect -1025 -288 -991 288
rect -929 -288 -895 288
rect -833 -288 -799 288
rect -737 -288 -703 288
rect -641 -288 -607 288
rect -545 -288 -511 288
rect -449 -288 -415 288
rect -353 -288 -319 288
rect -257 -288 -223 288
rect -161 -288 -127 288
rect -65 -288 -31 288
rect 31 -288 65 288
rect 127 -288 161 288
rect 223 -288 257 288
rect 319 -288 353 288
rect 415 -288 449 288
rect 511 -288 545 288
rect 607 -288 641 288
rect 703 -288 737 288
rect 799 -288 833 288
rect 895 -288 929 288
rect 991 -288 1025 288
rect 1087 -288 1121 288
rect 1183 -288 1217 288
rect 1279 -288 1313 288
rect -875 -395 875 -360
<< metal1 >>
rect -1280 395 -930 415
rect -1280 360 -1260 395
rect -950 360 -930 395
rect -1280 340 -930 360
rect 930 395 1280 415
rect 930 360 950 395
rect 1260 360 1280 395
rect 930 340 1280 360
rect -1319 288 -1273 300
rect -1319 -288 -1313 288
rect -1279 -288 -1273 288
rect -1319 -300 -1273 -288
rect -1223 288 -1177 300
rect -1223 -288 -1217 288
rect -1183 -288 -1177 288
rect -1223 -300 -1177 -288
rect -1127 288 -1081 300
rect -1127 -288 -1121 288
rect -1087 -288 -1081 288
rect -1127 -300 -1081 -288
rect -1031 288 -985 300
rect -1031 -288 -1025 288
rect -991 -288 -985 288
rect -1031 -300 -985 -288
rect -935 288 -889 300
rect -935 -288 -929 288
rect -895 -288 -889 288
rect -935 -300 -889 -288
rect -839 288 -793 300
rect -839 -288 -833 288
rect -799 -288 -793 288
rect -839 -300 -793 -288
rect -743 288 -697 300
rect -743 -288 -737 288
rect -703 -288 -697 288
rect -743 -300 -697 -288
rect -647 288 -601 300
rect -647 -288 -641 288
rect -607 -288 -601 288
rect -647 -300 -601 -288
rect -551 288 -505 300
rect -551 -288 -545 288
rect -511 -288 -505 288
rect -551 -300 -505 -288
rect -455 288 -409 300
rect -455 -288 -449 288
rect -415 -288 -409 288
rect -455 -300 -409 -288
rect -359 288 -313 300
rect -359 -288 -353 288
rect -319 -288 -313 288
rect -359 -300 -313 -288
rect -263 288 -217 300
rect -263 -288 -257 288
rect -223 -288 -217 288
rect -263 -300 -217 -288
rect -167 288 -121 300
rect -167 -288 -161 288
rect -127 -288 -121 288
rect -167 -300 -121 -288
rect -71 288 -25 300
rect -71 -288 -65 288
rect -31 -288 -25 288
rect -71 -300 -25 -288
rect 25 288 71 300
rect 25 -288 31 288
rect 65 -288 71 288
rect 25 -300 71 -288
rect 121 288 167 300
rect 121 -288 127 288
rect 161 -288 167 288
rect 121 -300 167 -288
rect 217 288 263 300
rect 217 -288 223 288
rect 257 -288 263 288
rect 217 -300 263 -288
rect 313 288 359 300
rect 313 -288 319 288
rect 353 -288 359 288
rect 313 -300 359 -288
rect 409 288 455 300
rect 409 -288 415 288
rect 449 -288 455 288
rect 409 -300 455 -288
rect 505 288 551 300
rect 505 -288 511 288
rect 545 -288 551 288
rect 505 -300 551 -288
rect 601 288 647 300
rect 601 -288 607 288
rect 641 -288 647 288
rect 601 -300 647 -288
rect 697 288 743 300
rect 697 -288 703 288
rect 737 -288 743 288
rect 697 -300 743 -288
rect 793 288 839 300
rect 793 -288 799 288
rect 833 -288 839 288
rect 793 -300 839 -288
rect 889 288 935 300
rect 889 -288 895 288
rect 929 -288 935 288
rect 889 -300 935 -288
rect 985 288 1031 300
rect 985 -288 991 288
rect 1025 -288 1031 288
rect 985 -300 1031 -288
rect 1081 288 1127 300
rect 1081 -288 1087 288
rect 1121 -288 1127 288
rect 1081 -300 1127 -288
rect 1177 288 1223 300
rect 1177 -288 1183 288
rect 1217 -288 1223 288
rect 1177 -300 1223 -288
rect 1273 288 1319 300
rect 1273 -288 1279 288
rect 1313 -288 1319 288
rect 1273 -300 1319 -288
rect -895 -360 895 -340
rect -895 -395 -875 -360
rect 875 -395 895 -360
rect -895 -415 895 -395
<< labels >>
rlabel nsubdiffcont 0 -466 0 -466 0 B
port 1 nsew
rlabel pdiffc -1296 0 -1296 0 0 D0
port 2 nsew
rlabel pdiffc -1200 0 -1200 0 0 S1
port 4 nsew
rlabel pdiffc -1104 0 -1104 0 0 D2
port 6 nsew
rlabel pdiffc -1008 0 -1008 0 0 S3
port 8 nsew
rlabel pdiffc -912 0 -912 0 0 D4
port 10 nsew
rlabel polycont -864 -364 -864 -364 0 G4
port 11 nsew
rlabel pdiffc -816 0 -816 0 0 S5
port 12 nsew
rlabel pdiffc -720 0 -720 0 0 D6
port 14 nsew
rlabel polycont -672 -364 -672 -364 0 G6
port 15 nsew
rlabel pdiffc -624 0 -624 0 0 S7
port 16 nsew
rlabel pdiffc -528 0 -528 0 0 D8
port 18 nsew
rlabel polycont -480 -364 -480 -364 0 G8
port 19 nsew
rlabel pdiffc -432 0 -432 0 0 S9
port 20 nsew
rlabel pdiffc -336 0 -336 0 0 D10
port 22 nsew
rlabel polycont -288 -364 -288 -364 0 G10
port 23 nsew
rlabel pdiffc -240 0 -240 0 0 S11
port 24 nsew
rlabel pdiffc -144 0 -144 0 0 D12
port 26 nsew
rlabel polycont -96 -364 -96 -364 0 G12
port 27 nsew
rlabel pdiffc -48 0 -48 0 0 S13
port 28 nsew
rlabel pdiffc 48 0 48 0 0 D14
port 30 nsew
rlabel polycont 96 -364 96 -364 0 G14
port 31 nsew
rlabel pdiffc 144 0 144 0 0 S15
port 32 nsew
rlabel pdiffc 240 0 240 0 0 D16
port 34 nsew
rlabel polycont 288 -364 288 -364 0 G16
port 35 nsew
rlabel pdiffc 336 0 336 0 0 S17
port 36 nsew
rlabel pdiffc 432 0 432 0 0 D18
port 38 nsew
rlabel polycont 480 -364 480 -364 0 G18
port 39 nsew
rlabel pdiffc 528 0 528 0 0 S19
port 40 nsew
rlabel pdiffc 624 0 624 0 0 D20
port 42 nsew
rlabel polycont 672 -364 672 -364 0 G20
port 43 nsew
rlabel pdiffc 720 0 720 0 0 S21
port 44 nsew
rlabel pdiffc 816 0 816 0 0 D22
port 46 nsew
rlabel polycont 864 -364 864 -364 0 G22
port 47 nsew
rlabel pdiffc 912 0 912 0 0 S23
port 48 nsew
rlabel polycont 960 364 960 364 0 G23
port 49 nsew
rlabel pdiffc 1008 0 1008 0 0 D24
port 50 nsew
rlabel pdiffc 1104 0 1104 0 0 S25
port 52 nsew
rlabel polycont 1152 364 1152 364 0 G25
port 53 nsew
rlabel pdiffc 1200 0 1200 0 0 D26
port 54 nsew
rlabel pdiffc 1296 0 1296 0 0 S26
port 55 nsew
<< properties >>
string FIXED_BBOX -1410 -466 1410 466
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3 l 0.15 m 1 nf 27 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
