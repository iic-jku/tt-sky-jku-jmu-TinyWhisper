magic
tech sky130A
magscale 1 2
timestamp 1762641840
<< pwell >>
rect -941 -510 941 510
<< nmoslvt >>
rect -745 -300 -545 300
rect -487 -300 -287 300
rect -229 -300 -29 300
rect 29 -300 229 300
rect 287 -300 487 300
rect 545 -300 745 300
<< ndiff >>
rect -803 288 -745 300
rect -803 -288 -791 288
rect -757 -288 -745 288
rect -803 -300 -745 -288
rect -545 288 -487 300
rect -545 -288 -533 288
rect -499 -288 -487 288
rect -545 -300 -487 -288
rect -287 288 -229 300
rect -287 -288 -275 288
rect -241 -288 -229 288
rect -287 -300 -229 -288
rect -29 288 29 300
rect -29 -288 -17 288
rect 17 -288 29 288
rect -29 -300 29 -288
rect 229 288 287 300
rect 229 -288 241 288
rect 275 -288 287 288
rect 229 -300 287 -288
rect 487 288 545 300
rect 487 -288 499 288
rect 533 -288 545 288
rect 487 -300 545 -288
rect 745 288 803 300
rect 745 -288 757 288
rect 791 -288 803 288
rect 745 -300 803 -288
<< ndiffc >>
rect -791 -288 -757 288
rect -533 -288 -499 288
rect -275 -288 -241 288
rect -17 -288 17 288
rect 241 -288 275 288
rect 499 -288 533 288
rect 757 -288 791 288
<< psubdiff >>
rect -905 440 -809 474
rect 809 440 905 474
rect -905 378 -871 440
rect 871 378 905 440
rect -905 -440 -871 -378
rect 871 -440 905 -378
rect -905 -474 -809 -440
rect 809 -474 905 -440
<< psubdiffcont >>
rect -809 440 809 474
rect -905 -378 -871 378
rect 871 -378 905 378
rect -809 -474 809 -440
<< poly >>
rect -487 372 -287 388
rect -487 338 -471 372
rect -303 338 -287 372
rect -745 300 -545 335
rect -487 300 -287 338
rect -229 372 -29 388
rect -229 338 -213 372
rect -45 338 -29 372
rect -229 300 -29 338
rect 29 372 229 388
rect 29 338 45 372
rect 213 338 229 372
rect 29 300 229 338
rect 287 372 487 388
rect 287 338 303 372
rect 471 338 487 372
rect 287 300 487 338
rect 545 300 745 335
rect -745 -338 -545 -300
rect -487 -335 -287 -300
rect -229 -335 -29 -300
rect 29 -335 229 -300
rect 287 -335 487 -300
rect -745 -372 -729 -338
rect -561 -372 -545 -338
rect -745 -388 -545 -372
rect 545 -338 745 -300
rect 545 -372 561 -338
rect 729 -372 745 -338
rect 545 -388 745 -372
<< polycont >>
rect -471 338 -303 372
rect -213 338 -45 372
rect 45 338 213 372
rect 303 338 471 372
rect -729 -372 -561 -338
rect 561 -372 729 -338
<< locali >>
rect -905 440 -809 474
rect 809 440 905 474
rect -905 378 -871 440
rect 871 378 905 440
rect -487 338 -471 372
rect -303 338 -287 372
rect -229 338 -213 372
rect -45 338 -29 372
rect 29 338 45 372
rect 213 338 229 372
rect 287 338 303 372
rect 471 338 487 372
rect -791 288 -757 304
rect -791 -304 -757 -288
rect -533 288 -499 304
rect -533 -304 -499 -288
rect -275 288 -241 304
rect -275 -304 -241 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 241 288 275 304
rect 241 -304 275 -288
rect 499 288 533 304
rect 499 -304 533 -288
rect 757 288 791 304
rect 757 -304 791 -288
rect -745 -372 -729 -338
rect -561 -372 -545 -338
rect 545 -372 561 -338
rect 729 -372 745 -338
rect -905 -440 -871 -378
rect 871 -440 905 -378
rect -905 -474 -809 -440
rect 809 -474 905 -440
<< viali >>
rect -471 338 -303 372
rect -213 338 -45 372
rect 45 338 213 372
rect 303 338 471 372
rect -791 -288 -757 288
rect -533 -288 -499 288
rect -275 -288 -241 288
rect -17 -288 17 288
rect 241 -288 275 288
rect 499 -288 533 288
rect 757 -288 791 288
rect -729 -372 -561 -338
rect 561 -372 729 -338
<< metal1 >>
rect -483 372 -291 378
rect -483 338 -471 372
rect -303 338 -291 372
rect -483 332 -291 338
rect -225 372 -33 378
rect -225 338 -213 372
rect -45 338 -33 372
rect -225 332 -33 338
rect 33 372 225 378
rect 33 338 45 372
rect 213 338 225 372
rect 33 332 225 338
rect 291 372 483 378
rect 291 338 303 372
rect 471 338 483 372
rect 291 332 483 338
rect -797 288 -751 300
rect -797 -288 -791 288
rect -757 -288 -751 288
rect -797 -300 -751 -288
rect -539 288 -493 300
rect -539 -288 -533 288
rect -499 -288 -493 288
rect -539 -300 -493 -288
rect -281 288 -235 300
rect -281 -288 -275 288
rect -241 -288 -235 288
rect -281 -300 -235 -288
rect -23 288 23 300
rect -23 -288 -17 288
rect 17 -288 23 288
rect -23 -300 23 -288
rect 235 288 281 300
rect 235 -288 241 288
rect 275 -288 281 288
rect 235 -300 281 -288
rect 493 288 539 300
rect 493 -288 499 288
rect 533 -288 539 288
rect 493 -300 539 -288
rect 751 288 797 300
rect 751 -288 757 288
rect 791 -288 797 288
rect 751 -300 797 -288
rect -741 -338 -549 -332
rect -741 -372 -729 -338
rect -561 -372 -549 -338
rect -741 -378 -549 -372
rect 549 -338 741 -332
rect 549 -372 561 -338
rect 729 -372 741 -338
rect 549 -378 741 -372
<< labels >>
rlabel psubdiffcont 0 -457 0 -457 0 B
port 1 nsew
rlabel ndiffc -774 0 -774 0 0 D0
port 2 nsew
rlabel ndiffc -516 0 -516 0 0 S1
port 4 nsew
rlabel polycont -387 355 -387 355 0 G1
port 5 nsew
rlabel ndiffc -258 0 -258 0 0 D2
port 6 nsew
rlabel polycont -129 355 -129 355 0 G2
port 7 nsew
rlabel ndiffc 0 0 0 0 0 S3
port 8 nsew
rlabel polycont 129 355 129 355 0 G3
port 9 nsew
rlabel ndiffc 258 0 258 0 0 D4
port 10 nsew
rlabel polycont 387 355 387 355 0 G4
port 11 nsew
rlabel ndiffc 516 0 516 0 0 S5
port 12 nsew
<< properties >>
string FIXED_BBOX -888 -457 888 457
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 3 l 1 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
