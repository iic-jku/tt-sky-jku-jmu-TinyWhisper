magic
tech sky130A
magscale 1 2
timestamp 1762706219
<< metal3 >>
rect -516 2312 516 2340
rect -516 1688 432 2312
rect 496 1688 516 2312
rect -516 1660 516 1688
rect -516 1312 516 1340
rect -516 688 432 1312
rect 496 688 516 1312
rect -516 660 516 688
rect -516 312 516 340
rect -516 -312 432 312
rect 496 -312 516 312
rect -516 -340 516 -312
rect -516 -688 516 -660
rect -516 -1312 432 -688
rect 496 -1312 516 -688
rect -516 -1340 516 -1312
rect -516 -1688 516 -1660
rect -516 -2312 432 -1688
rect 496 -2312 516 -1688
rect -516 -2340 516 -2312
<< via3 >>
rect 432 1688 496 2312
rect 432 688 496 1312
rect 432 -312 496 312
rect 432 -1312 496 -688
rect 432 -2312 496 -1688
<< mimcap >>
rect -476 2260 124 2300
rect -476 1740 -436 2260
rect 84 1740 124 2260
rect -476 1700 124 1740
rect -476 1260 124 1300
rect -476 740 -436 1260
rect 84 740 124 1260
rect -476 700 124 740
rect -476 260 124 300
rect -476 -260 -436 260
rect 84 -260 124 260
rect -476 -300 124 -260
rect -476 -740 124 -700
rect -476 -1260 -436 -740
rect 84 -1260 124 -740
rect -476 -1300 124 -1260
rect -476 -1740 124 -1700
rect -476 -2260 -436 -1740
rect 84 -2260 124 -1740
rect -476 -2300 124 -2260
<< mimcapcontact >>
rect -436 1740 84 2260
rect -436 740 84 1260
rect -436 -260 84 260
rect -436 -1260 84 -740
rect -436 -2260 84 -1740
<< metal4 >>
rect -228 2261 -124 2500
rect 412 2312 516 2500
rect -437 2260 85 2261
rect -437 1740 -436 2260
rect 84 1740 85 2260
rect -437 1739 85 1740
rect -228 1261 -124 1739
rect 412 1688 432 2312
rect 496 1688 516 2312
rect 412 1312 516 1688
rect -437 1260 85 1261
rect -437 740 -436 1260
rect 84 740 85 1260
rect -437 739 85 740
rect -228 261 -124 739
rect 412 688 432 1312
rect 496 688 516 1312
rect 412 312 516 688
rect -437 260 85 261
rect -437 -260 -436 260
rect 84 -260 85 260
rect -437 -261 85 -260
rect -228 -739 -124 -261
rect 412 -312 432 312
rect 496 -312 516 312
rect 412 -688 516 -312
rect -437 -740 85 -739
rect -437 -1260 -436 -740
rect 84 -1260 85 -740
rect -437 -1261 85 -1260
rect -228 -1739 -124 -1261
rect 412 -1312 432 -688
rect 496 -1312 516 -688
rect 412 -1688 516 -1312
rect -437 -1740 85 -1739
rect -437 -2260 -436 -1740
rect 84 -2260 85 -1740
rect -437 -2261 85 -2260
rect -228 -2500 -124 -2261
rect 412 -2312 432 -1688
rect 496 -2312 516 -1688
rect 412 -2500 516 -2312
<< labels >>
rlabel via3 464 -2000 464 -2000 0 C2
port 1 nsew
rlabel mimcapcontact -176 -2000 -176 -2000 0 C1
port 2 nsew
<< properties >>
string FIXED_BBOX -516 1660 164 2340
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 3.00 l 3.00 val 20.28 carea 2.00 cperi 0.19 class capacitor nx 1 ny 5 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100 stack 1 doports 1
<< end >>
