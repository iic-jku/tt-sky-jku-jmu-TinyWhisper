magic
tech sky130A
magscale 1 2
timestamp 1762702375
<< metal3 >>
rect -11553 1812 -10521 1840
rect -11553 1188 -10605 1812
rect -10541 1188 -10521 1812
rect -11553 1160 -10521 1188
rect -9855 1812 -8823 1840
rect -9855 1188 -8907 1812
rect -8843 1188 -8823 1812
rect -9855 1160 -8823 1188
rect -8157 1812 -7125 1840
rect -8157 1188 -7209 1812
rect -7145 1188 -7125 1812
rect -8157 1160 -7125 1188
rect -6459 1812 -5427 1840
rect -6459 1188 -5511 1812
rect -5447 1188 -5427 1812
rect -6459 1160 -5427 1188
rect -4761 1812 -3729 1840
rect -4761 1188 -3813 1812
rect -3749 1188 -3729 1812
rect -4761 1160 -3729 1188
rect -3063 1812 -2031 1840
rect -3063 1188 -2115 1812
rect -2051 1188 -2031 1812
rect -3063 1160 -2031 1188
rect -1365 1812 -333 1840
rect -1365 1188 -417 1812
rect -353 1188 -333 1812
rect -1365 1160 -333 1188
rect 333 1812 1365 1840
rect 333 1188 1281 1812
rect 1345 1188 1365 1812
rect 333 1160 1365 1188
rect 2031 1812 3063 1840
rect 2031 1188 2979 1812
rect 3043 1188 3063 1812
rect 2031 1160 3063 1188
rect 3729 1812 4761 1840
rect 3729 1188 4677 1812
rect 4741 1188 4761 1812
rect 3729 1160 4761 1188
rect 5427 1812 6459 1840
rect 5427 1188 6375 1812
rect 6439 1188 6459 1812
rect 5427 1160 6459 1188
rect 7125 1812 8157 1840
rect 7125 1188 8073 1812
rect 8137 1188 8157 1812
rect 7125 1160 8157 1188
rect 8823 1812 9855 1840
rect 8823 1188 9771 1812
rect 9835 1188 9855 1812
rect 8823 1160 9855 1188
rect 10521 1812 11553 1840
rect 10521 1188 11469 1812
rect 11533 1188 11553 1812
rect 10521 1160 11553 1188
rect -11553 812 -10521 840
rect -11553 188 -10605 812
rect -10541 188 -10521 812
rect -11553 160 -10521 188
rect -9855 812 -8823 840
rect -9855 188 -8907 812
rect -8843 188 -8823 812
rect -9855 160 -8823 188
rect -8157 812 -7125 840
rect -8157 188 -7209 812
rect -7145 188 -7125 812
rect -8157 160 -7125 188
rect -6459 812 -5427 840
rect -6459 188 -5511 812
rect -5447 188 -5427 812
rect -6459 160 -5427 188
rect -4761 812 -3729 840
rect -4761 188 -3813 812
rect -3749 188 -3729 812
rect -4761 160 -3729 188
rect -3063 812 -2031 840
rect -3063 188 -2115 812
rect -2051 188 -2031 812
rect -3063 160 -2031 188
rect -1365 812 -333 840
rect -1365 188 -417 812
rect -353 188 -333 812
rect -1365 160 -333 188
rect 333 812 1365 840
rect 333 188 1281 812
rect 1345 188 1365 812
rect 333 160 1365 188
rect 2031 812 3063 840
rect 2031 188 2979 812
rect 3043 188 3063 812
rect 2031 160 3063 188
rect 3729 812 4761 840
rect 3729 188 4677 812
rect 4741 188 4761 812
rect 3729 160 4761 188
rect 5427 812 6459 840
rect 5427 188 6375 812
rect 6439 188 6459 812
rect 5427 160 6459 188
rect 7125 812 8157 840
rect 7125 188 8073 812
rect 8137 188 8157 812
rect 7125 160 8157 188
rect 8823 812 9855 840
rect 8823 188 9771 812
rect 9835 188 9855 812
rect 8823 160 9855 188
rect 10521 812 11553 840
rect 10521 188 11469 812
rect 11533 188 11553 812
rect 10521 160 11553 188
rect -11553 -188 -10521 -160
rect -11553 -812 -10605 -188
rect -10541 -812 -10521 -188
rect -11553 -840 -10521 -812
rect -9855 -188 -8823 -160
rect -9855 -812 -8907 -188
rect -8843 -812 -8823 -188
rect -9855 -840 -8823 -812
rect -8157 -188 -7125 -160
rect -8157 -812 -7209 -188
rect -7145 -812 -7125 -188
rect -8157 -840 -7125 -812
rect -6459 -188 -5427 -160
rect -6459 -812 -5511 -188
rect -5447 -812 -5427 -188
rect -6459 -840 -5427 -812
rect -4761 -188 -3729 -160
rect -4761 -812 -3813 -188
rect -3749 -812 -3729 -188
rect -4761 -840 -3729 -812
rect -3063 -188 -2031 -160
rect -3063 -812 -2115 -188
rect -2051 -812 -2031 -188
rect -3063 -840 -2031 -812
rect -1365 -188 -333 -160
rect -1365 -812 -417 -188
rect -353 -812 -333 -188
rect -1365 -840 -333 -812
rect 333 -188 1365 -160
rect 333 -812 1281 -188
rect 1345 -812 1365 -188
rect 333 -840 1365 -812
rect 2031 -188 3063 -160
rect 2031 -812 2979 -188
rect 3043 -812 3063 -188
rect 2031 -840 3063 -812
rect 3729 -188 4761 -160
rect 3729 -812 4677 -188
rect 4741 -812 4761 -188
rect 3729 -840 4761 -812
rect 5427 -188 6459 -160
rect 5427 -812 6375 -188
rect 6439 -812 6459 -188
rect 5427 -840 6459 -812
rect 7125 -188 8157 -160
rect 7125 -812 8073 -188
rect 8137 -812 8157 -188
rect 7125 -840 8157 -812
rect 8823 -188 9855 -160
rect 8823 -812 9771 -188
rect 9835 -812 9855 -188
rect 8823 -840 9855 -812
rect 10521 -188 11553 -160
rect 10521 -812 11469 -188
rect 11533 -812 11553 -188
rect 10521 -840 11553 -812
rect -11553 -1188 -10521 -1160
rect -11553 -1812 -10605 -1188
rect -10541 -1812 -10521 -1188
rect -11553 -1840 -10521 -1812
rect -9855 -1188 -8823 -1160
rect -9855 -1812 -8907 -1188
rect -8843 -1812 -8823 -1188
rect -9855 -1840 -8823 -1812
rect -8157 -1188 -7125 -1160
rect -8157 -1812 -7209 -1188
rect -7145 -1812 -7125 -1188
rect -8157 -1840 -7125 -1812
rect -6459 -1188 -5427 -1160
rect -6459 -1812 -5511 -1188
rect -5447 -1812 -5427 -1188
rect -6459 -1840 -5427 -1812
rect -4761 -1188 -3729 -1160
rect -4761 -1812 -3813 -1188
rect -3749 -1812 -3729 -1188
rect -4761 -1840 -3729 -1812
rect -3063 -1188 -2031 -1160
rect -3063 -1812 -2115 -1188
rect -2051 -1812 -2031 -1188
rect -3063 -1840 -2031 -1812
rect -1365 -1188 -333 -1160
rect -1365 -1812 -417 -1188
rect -353 -1812 -333 -1188
rect -1365 -1840 -333 -1812
rect 333 -1188 1365 -1160
rect 333 -1812 1281 -1188
rect 1345 -1812 1365 -1188
rect 333 -1840 1365 -1812
rect 2031 -1188 3063 -1160
rect 2031 -1812 2979 -1188
rect 3043 -1812 3063 -1188
rect 2031 -1840 3063 -1812
rect 3729 -1188 4761 -1160
rect 3729 -1812 4677 -1188
rect 4741 -1812 4761 -1188
rect 3729 -1840 4761 -1812
rect 5427 -1188 6459 -1160
rect 5427 -1812 6375 -1188
rect 6439 -1812 6459 -1188
rect 5427 -1840 6459 -1812
rect 7125 -1188 8157 -1160
rect 7125 -1812 8073 -1188
rect 8137 -1812 8157 -1188
rect 7125 -1840 8157 -1812
rect 8823 -1188 9855 -1160
rect 8823 -1812 9771 -1188
rect 9835 -1812 9855 -1188
rect 8823 -1840 9855 -1812
rect 10521 -1188 11553 -1160
rect 10521 -1812 11469 -1188
rect 11533 -1812 11553 -1188
rect 10521 -1840 11553 -1812
<< via3 >>
rect -10605 1188 -10541 1812
rect -8907 1188 -8843 1812
rect -7209 1188 -7145 1812
rect -5511 1188 -5447 1812
rect -3813 1188 -3749 1812
rect -2115 1188 -2051 1812
rect -417 1188 -353 1812
rect 1281 1188 1345 1812
rect 2979 1188 3043 1812
rect 4677 1188 4741 1812
rect 6375 1188 6439 1812
rect 8073 1188 8137 1812
rect 9771 1188 9835 1812
rect 11469 1188 11533 1812
rect -10605 188 -10541 812
rect -8907 188 -8843 812
rect -7209 188 -7145 812
rect -5511 188 -5447 812
rect -3813 188 -3749 812
rect -2115 188 -2051 812
rect -417 188 -353 812
rect 1281 188 1345 812
rect 2979 188 3043 812
rect 4677 188 4741 812
rect 6375 188 6439 812
rect 8073 188 8137 812
rect 9771 188 9835 812
rect 11469 188 11533 812
rect -10605 -812 -10541 -188
rect -8907 -812 -8843 -188
rect -7209 -812 -7145 -188
rect -5511 -812 -5447 -188
rect -3813 -812 -3749 -188
rect -2115 -812 -2051 -188
rect -417 -812 -353 -188
rect 1281 -812 1345 -188
rect 2979 -812 3043 -188
rect 4677 -812 4741 -188
rect 6375 -812 6439 -188
rect 8073 -812 8137 -188
rect 9771 -812 9835 -188
rect 11469 -812 11533 -188
rect -10605 -1812 -10541 -1188
rect -8907 -1812 -8843 -1188
rect -7209 -1812 -7145 -1188
rect -5511 -1812 -5447 -1188
rect -3813 -1812 -3749 -1188
rect -2115 -1812 -2051 -1188
rect -417 -1812 -353 -1188
rect 1281 -1812 1345 -1188
rect 2979 -1812 3043 -1188
rect 4677 -1812 4741 -1188
rect 6375 -1812 6439 -1188
rect 8073 -1812 8137 -1188
rect 9771 -1812 9835 -1188
rect 11469 -1812 11533 -1188
<< mimcap >>
rect -11513 1760 -10913 1800
rect -11513 1240 -11473 1760
rect -10953 1240 -10913 1760
rect -11513 1200 -10913 1240
rect -9815 1760 -9215 1800
rect -9815 1240 -9775 1760
rect -9255 1240 -9215 1760
rect -9815 1200 -9215 1240
rect -8117 1760 -7517 1800
rect -8117 1240 -8077 1760
rect -7557 1240 -7517 1760
rect -8117 1200 -7517 1240
rect -6419 1760 -5819 1800
rect -6419 1240 -6379 1760
rect -5859 1240 -5819 1760
rect -6419 1200 -5819 1240
rect -4721 1760 -4121 1800
rect -4721 1240 -4681 1760
rect -4161 1240 -4121 1760
rect -4721 1200 -4121 1240
rect -3023 1760 -2423 1800
rect -3023 1240 -2983 1760
rect -2463 1240 -2423 1760
rect -3023 1200 -2423 1240
rect -1325 1760 -725 1800
rect -1325 1240 -1285 1760
rect -765 1240 -725 1760
rect -1325 1200 -725 1240
rect 373 1760 973 1800
rect 373 1240 413 1760
rect 933 1240 973 1760
rect 373 1200 973 1240
rect 2071 1760 2671 1800
rect 2071 1240 2111 1760
rect 2631 1240 2671 1760
rect 2071 1200 2671 1240
rect 3769 1760 4369 1800
rect 3769 1240 3809 1760
rect 4329 1240 4369 1760
rect 3769 1200 4369 1240
rect 5467 1760 6067 1800
rect 5467 1240 5507 1760
rect 6027 1240 6067 1760
rect 5467 1200 6067 1240
rect 7165 1760 7765 1800
rect 7165 1240 7205 1760
rect 7725 1240 7765 1760
rect 7165 1200 7765 1240
rect 8863 1760 9463 1800
rect 8863 1240 8903 1760
rect 9423 1240 9463 1760
rect 8863 1200 9463 1240
rect 10561 1760 11161 1800
rect 10561 1240 10601 1760
rect 11121 1240 11161 1760
rect 10561 1200 11161 1240
rect -11513 760 -10913 800
rect -11513 240 -11473 760
rect -10953 240 -10913 760
rect -11513 200 -10913 240
rect -9815 760 -9215 800
rect -9815 240 -9775 760
rect -9255 240 -9215 760
rect -9815 200 -9215 240
rect -8117 760 -7517 800
rect -8117 240 -8077 760
rect -7557 240 -7517 760
rect -8117 200 -7517 240
rect -6419 760 -5819 800
rect -6419 240 -6379 760
rect -5859 240 -5819 760
rect -6419 200 -5819 240
rect -4721 760 -4121 800
rect -4721 240 -4681 760
rect -4161 240 -4121 760
rect -4721 200 -4121 240
rect -3023 760 -2423 800
rect -3023 240 -2983 760
rect -2463 240 -2423 760
rect -3023 200 -2423 240
rect -1325 760 -725 800
rect -1325 240 -1285 760
rect -765 240 -725 760
rect -1325 200 -725 240
rect 373 760 973 800
rect 373 240 413 760
rect 933 240 973 760
rect 373 200 973 240
rect 2071 760 2671 800
rect 2071 240 2111 760
rect 2631 240 2671 760
rect 2071 200 2671 240
rect 3769 760 4369 800
rect 3769 240 3809 760
rect 4329 240 4369 760
rect 3769 200 4369 240
rect 5467 760 6067 800
rect 5467 240 5507 760
rect 6027 240 6067 760
rect 5467 200 6067 240
rect 7165 760 7765 800
rect 7165 240 7205 760
rect 7725 240 7765 760
rect 7165 200 7765 240
rect 8863 760 9463 800
rect 8863 240 8903 760
rect 9423 240 9463 760
rect 8863 200 9463 240
rect 10561 760 11161 800
rect 10561 240 10601 760
rect 11121 240 11161 760
rect 10561 200 11161 240
rect -11513 -240 -10913 -200
rect -11513 -760 -11473 -240
rect -10953 -760 -10913 -240
rect -11513 -800 -10913 -760
rect -9815 -240 -9215 -200
rect -9815 -760 -9775 -240
rect -9255 -760 -9215 -240
rect -9815 -800 -9215 -760
rect -8117 -240 -7517 -200
rect -8117 -760 -8077 -240
rect -7557 -760 -7517 -240
rect -8117 -800 -7517 -760
rect -6419 -240 -5819 -200
rect -6419 -760 -6379 -240
rect -5859 -760 -5819 -240
rect -6419 -800 -5819 -760
rect -4721 -240 -4121 -200
rect -4721 -760 -4681 -240
rect -4161 -760 -4121 -240
rect -4721 -800 -4121 -760
rect -3023 -240 -2423 -200
rect -3023 -760 -2983 -240
rect -2463 -760 -2423 -240
rect -3023 -800 -2423 -760
rect -1325 -240 -725 -200
rect -1325 -760 -1285 -240
rect -765 -760 -725 -240
rect -1325 -800 -725 -760
rect 373 -240 973 -200
rect 373 -760 413 -240
rect 933 -760 973 -240
rect 373 -800 973 -760
rect 2071 -240 2671 -200
rect 2071 -760 2111 -240
rect 2631 -760 2671 -240
rect 2071 -800 2671 -760
rect 3769 -240 4369 -200
rect 3769 -760 3809 -240
rect 4329 -760 4369 -240
rect 3769 -800 4369 -760
rect 5467 -240 6067 -200
rect 5467 -760 5507 -240
rect 6027 -760 6067 -240
rect 5467 -800 6067 -760
rect 7165 -240 7765 -200
rect 7165 -760 7205 -240
rect 7725 -760 7765 -240
rect 7165 -800 7765 -760
rect 8863 -240 9463 -200
rect 8863 -760 8903 -240
rect 9423 -760 9463 -240
rect 8863 -800 9463 -760
rect 10561 -240 11161 -200
rect 10561 -760 10601 -240
rect 11121 -760 11161 -240
rect 10561 -800 11161 -760
rect -11513 -1240 -10913 -1200
rect -11513 -1760 -11473 -1240
rect -10953 -1760 -10913 -1240
rect -11513 -1800 -10913 -1760
rect -9815 -1240 -9215 -1200
rect -9815 -1760 -9775 -1240
rect -9255 -1760 -9215 -1240
rect -9815 -1800 -9215 -1760
rect -8117 -1240 -7517 -1200
rect -8117 -1760 -8077 -1240
rect -7557 -1760 -7517 -1240
rect -8117 -1800 -7517 -1760
rect -6419 -1240 -5819 -1200
rect -6419 -1760 -6379 -1240
rect -5859 -1760 -5819 -1240
rect -6419 -1800 -5819 -1760
rect -4721 -1240 -4121 -1200
rect -4721 -1760 -4681 -1240
rect -4161 -1760 -4121 -1240
rect -4721 -1800 -4121 -1760
rect -3023 -1240 -2423 -1200
rect -3023 -1760 -2983 -1240
rect -2463 -1760 -2423 -1240
rect -3023 -1800 -2423 -1760
rect -1325 -1240 -725 -1200
rect -1325 -1760 -1285 -1240
rect -765 -1760 -725 -1240
rect -1325 -1800 -725 -1760
rect 373 -1240 973 -1200
rect 373 -1760 413 -1240
rect 933 -1760 973 -1240
rect 373 -1800 973 -1760
rect 2071 -1240 2671 -1200
rect 2071 -1760 2111 -1240
rect 2631 -1760 2671 -1240
rect 2071 -1800 2671 -1760
rect 3769 -1240 4369 -1200
rect 3769 -1760 3809 -1240
rect 4329 -1760 4369 -1240
rect 3769 -1800 4369 -1760
rect 5467 -1240 6067 -1200
rect 5467 -1760 5507 -1240
rect 6027 -1760 6067 -1240
rect 5467 -1800 6067 -1760
rect 7165 -1240 7765 -1200
rect 7165 -1760 7205 -1240
rect 7725 -1760 7765 -1240
rect 7165 -1800 7765 -1760
rect 8863 -1240 9463 -1200
rect 8863 -1760 8903 -1240
rect 9423 -1760 9463 -1240
rect 8863 -1800 9463 -1760
rect 10561 -1240 11161 -1200
rect 10561 -1760 10601 -1240
rect 11121 -1760 11161 -1240
rect 10561 -1800 11161 -1760
<< mimcapcontact >>
rect -11473 1240 -10953 1760
rect -9775 1240 -9255 1760
rect -8077 1240 -7557 1760
rect -6379 1240 -5859 1760
rect -4681 1240 -4161 1760
rect -2983 1240 -2463 1760
rect -1285 1240 -765 1760
rect 413 1240 933 1760
rect 2111 1240 2631 1760
rect 3809 1240 4329 1760
rect 5507 1240 6027 1760
rect 7205 1240 7725 1760
rect 8903 1240 9423 1760
rect 10601 1240 11121 1760
rect -11473 240 -10953 760
rect -9775 240 -9255 760
rect -8077 240 -7557 760
rect -6379 240 -5859 760
rect -4681 240 -4161 760
rect -2983 240 -2463 760
rect -1285 240 -765 760
rect 413 240 933 760
rect 2111 240 2631 760
rect 3809 240 4329 760
rect 5507 240 6027 760
rect 7205 240 7725 760
rect 8903 240 9423 760
rect 10601 240 11121 760
rect -11473 -760 -10953 -240
rect -9775 -760 -9255 -240
rect -8077 -760 -7557 -240
rect -6379 -760 -5859 -240
rect -4681 -760 -4161 -240
rect -2983 -760 -2463 -240
rect -1285 -760 -765 -240
rect 413 -760 933 -240
rect 2111 -760 2631 -240
rect 3809 -760 4329 -240
rect 5507 -760 6027 -240
rect 7205 -760 7725 -240
rect 8903 -760 9423 -240
rect 10601 -760 11121 -240
rect -11473 -1760 -10953 -1240
rect -9775 -1760 -9255 -1240
rect -8077 -1760 -7557 -1240
rect -6379 -1760 -5859 -1240
rect -4681 -1760 -4161 -1240
rect -2983 -1760 -2463 -1240
rect -1285 -1760 -765 -1240
rect 413 -1760 933 -1240
rect 2111 -1760 2631 -1240
rect 3809 -1760 4329 -1240
rect 5507 -1760 6027 -1240
rect 7205 -1760 7725 -1240
rect 8903 -1760 9423 -1240
rect 10601 -1760 11121 -1240
<< metal4 >>
rect -11265 1761 -11161 2000
rect -10625 1812 -10521 2000
rect -11474 1760 -10952 1761
rect -11474 1240 -11473 1760
rect -10953 1240 -10952 1760
rect -11474 1239 -10952 1240
rect -11265 761 -11161 1239
rect -10625 1188 -10605 1812
rect -10541 1188 -10521 1812
rect -9567 1761 -9463 2000
rect -8927 1812 -8823 2000
rect -9776 1760 -9254 1761
rect -9776 1240 -9775 1760
rect -9255 1240 -9254 1760
rect -9776 1239 -9254 1240
rect -10625 812 -10521 1188
rect -11474 760 -10952 761
rect -11474 240 -11473 760
rect -10953 240 -10952 760
rect -11474 239 -10952 240
rect -11265 -239 -11161 239
rect -10625 188 -10605 812
rect -10541 188 -10521 812
rect -9567 761 -9463 1239
rect -8927 1188 -8907 1812
rect -8843 1188 -8823 1812
rect -7869 1761 -7765 2000
rect -7229 1812 -7125 2000
rect -8078 1760 -7556 1761
rect -8078 1240 -8077 1760
rect -7557 1240 -7556 1760
rect -8078 1239 -7556 1240
rect -8927 812 -8823 1188
rect -9776 760 -9254 761
rect -9776 240 -9775 760
rect -9255 240 -9254 760
rect -9776 239 -9254 240
rect -10625 -188 -10521 188
rect -11474 -240 -10952 -239
rect -11474 -760 -11473 -240
rect -10953 -760 -10952 -240
rect -11474 -761 -10952 -760
rect -11265 -1239 -11161 -761
rect -10625 -812 -10605 -188
rect -10541 -812 -10521 -188
rect -9567 -239 -9463 239
rect -8927 188 -8907 812
rect -8843 188 -8823 812
rect -7869 761 -7765 1239
rect -7229 1188 -7209 1812
rect -7145 1188 -7125 1812
rect -6171 1761 -6067 2000
rect -5531 1812 -5427 2000
rect -6380 1760 -5858 1761
rect -6380 1240 -6379 1760
rect -5859 1240 -5858 1760
rect -6380 1239 -5858 1240
rect -7229 812 -7125 1188
rect -8078 760 -7556 761
rect -8078 240 -8077 760
rect -7557 240 -7556 760
rect -8078 239 -7556 240
rect -8927 -188 -8823 188
rect -9776 -240 -9254 -239
rect -9776 -760 -9775 -240
rect -9255 -760 -9254 -240
rect -9776 -761 -9254 -760
rect -10625 -1188 -10521 -812
rect -11474 -1240 -10952 -1239
rect -11474 -1760 -11473 -1240
rect -10953 -1760 -10952 -1240
rect -11474 -1761 -10952 -1760
rect -11265 -2000 -11161 -1761
rect -10625 -1812 -10605 -1188
rect -10541 -1812 -10521 -1188
rect -9567 -1239 -9463 -761
rect -8927 -812 -8907 -188
rect -8843 -812 -8823 -188
rect -7869 -239 -7765 239
rect -7229 188 -7209 812
rect -7145 188 -7125 812
rect -6171 761 -6067 1239
rect -5531 1188 -5511 1812
rect -5447 1188 -5427 1812
rect -4473 1761 -4369 2000
rect -3833 1812 -3729 2000
rect -4682 1760 -4160 1761
rect -4682 1240 -4681 1760
rect -4161 1240 -4160 1760
rect -4682 1239 -4160 1240
rect -5531 812 -5427 1188
rect -6380 760 -5858 761
rect -6380 240 -6379 760
rect -5859 240 -5858 760
rect -6380 239 -5858 240
rect -7229 -188 -7125 188
rect -8078 -240 -7556 -239
rect -8078 -760 -8077 -240
rect -7557 -760 -7556 -240
rect -8078 -761 -7556 -760
rect -8927 -1188 -8823 -812
rect -9776 -1240 -9254 -1239
rect -9776 -1760 -9775 -1240
rect -9255 -1760 -9254 -1240
rect -9776 -1761 -9254 -1760
rect -10625 -2000 -10521 -1812
rect -9567 -2000 -9463 -1761
rect -8927 -1812 -8907 -1188
rect -8843 -1812 -8823 -1188
rect -7869 -1239 -7765 -761
rect -7229 -812 -7209 -188
rect -7145 -812 -7125 -188
rect -6171 -239 -6067 239
rect -5531 188 -5511 812
rect -5447 188 -5427 812
rect -4473 761 -4369 1239
rect -3833 1188 -3813 1812
rect -3749 1188 -3729 1812
rect -2775 1761 -2671 2000
rect -2135 1812 -2031 2000
rect -2984 1760 -2462 1761
rect -2984 1240 -2983 1760
rect -2463 1240 -2462 1760
rect -2984 1239 -2462 1240
rect -3833 812 -3729 1188
rect -4682 760 -4160 761
rect -4682 240 -4681 760
rect -4161 240 -4160 760
rect -4682 239 -4160 240
rect -5531 -188 -5427 188
rect -6380 -240 -5858 -239
rect -6380 -760 -6379 -240
rect -5859 -760 -5858 -240
rect -6380 -761 -5858 -760
rect -7229 -1188 -7125 -812
rect -8078 -1240 -7556 -1239
rect -8078 -1760 -8077 -1240
rect -7557 -1760 -7556 -1240
rect -8078 -1761 -7556 -1760
rect -8927 -2000 -8823 -1812
rect -7869 -2000 -7765 -1761
rect -7229 -1812 -7209 -1188
rect -7145 -1812 -7125 -1188
rect -6171 -1239 -6067 -761
rect -5531 -812 -5511 -188
rect -5447 -812 -5427 -188
rect -4473 -239 -4369 239
rect -3833 188 -3813 812
rect -3749 188 -3729 812
rect -2775 761 -2671 1239
rect -2135 1188 -2115 1812
rect -2051 1188 -2031 1812
rect -1077 1761 -973 2000
rect -437 1812 -333 2000
rect -1286 1760 -764 1761
rect -1286 1240 -1285 1760
rect -765 1240 -764 1760
rect -1286 1239 -764 1240
rect -2135 812 -2031 1188
rect -2984 760 -2462 761
rect -2984 240 -2983 760
rect -2463 240 -2462 760
rect -2984 239 -2462 240
rect -3833 -188 -3729 188
rect -4682 -240 -4160 -239
rect -4682 -760 -4681 -240
rect -4161 -760 -4160 -240
rect -4682 -761 -4160 -760
rect -5531 -1188 -5427 -812
rect -6380 -1240 -5858 -1239
rect -6380 -1760 -6379 -1240
rect -5859 -1760 -5858 -1240
rect -6380 -1761 -5858 -1760
rect -7229 -2000 -7125 -1812
rect -6171 -2000 -6067 -1761
rect -5531 -1812 -5511 -1188
rect -5447 -1812 -5427 -1188
rect -4473 -1239 -4369 -761
rect -3833 -812 -3813 -188
rect -3749 -812 -3729 -188
rect -2775 -239 -2671 239
rect -2135 188 -2115 812
rect -2051 188 -2031 812
rect -1077 761 -973 1239
rect -437 1188 -417 1812
rect -353 1188 -333 1812
rect 621 1761 725 2000
rect 1261 1812 1365 2000
rect 412 1760 934 1761
rect 412 1240 413 1760
rect 933 1240 934 1760
rect 412 1239 934 1240
rect -437 812 -333 1188
rect -1286 760 -764 761
rect -1286 240 -1285 760
rect -765 240 -764 760
rect -1286 239 -764 240
rect -2135 -188 -2031 188
rect -2984 -240 -2462 -239
rect -2984 -760 -2983 -240
rect -2463 -760 -2462 -240
rect -2984 -761 -2462 -760
rect -3833 -1188 -3729 -812
rect -4682 -1240 -4160 -1239
rect -4682 -1760 -4681 -1240
rect -4161 -1760 -4160 -1240
rect -4682 -1761 -4160 -1760
rect -5531 -2000 -5427 -1812
rect -4473 -2000 -4369 -1761
rect -3833 -1812 -3813 -1188
rect -3749 -1812 -3729 -1188
rect -2775 -1239 -2671 -761
rect -2135 -812 -2115 -188
rect -2051 -812 -2031 -188
rect -1077 -239 -973 239
rect -437 188 -417 812
rect -353 188 -333 812
rect 621 761 725 1239
rect 1261 1188 1281 1812
rect 1345 1188 1365 1812
rect 2319 1761 2423 2000
rect 2959 1812 3063 2000
rect 2110 1760 2632 1761
rect 2110 1240 2111 1760
rect 2631 1240 2632 1760
rect 2110 1239 2632 1240
rect 1261 812 1365 1188
rect 412 760 934 761
rect 412 240 413 760
rect 933 240 934 760
rect 412 239 934 240
rect -437 -188 -333 188
rect -1286 -240 -764 -239
rect -1286 -760 -1285 -240
rect -765 -760 -764 -240
rect -1286 -761 -764 -760
rect -2135 -1188 -2031 -812
rect -2984 -1240 -2462 -1239
rect -2984 -1760 -2983 -1240
rect -2463 -1760 -2462 -1240
rect -2984 -1761 -2462 -1760
rect -3833 -2000 -3729 -1812
rect -2775 -2000 -2671 -1761
rect -2135 -1812 -2115 -1188
rect -2051 -1812 -2031 -1188
rect -1077 -1239 -973 -761
rect -437 -812 -417 -188
rect -353 -812 -333 -188
rect 621 -239 725 239
rect 1261 188 1281 812
rect 1345 188 1365 812
rect 2319 761 2423 1239
rect 2959 1188 2979 1812
rect 3043 1188 3063 1812
rect 4017 1761 4121 2000
rect 4657 1812 4761 2000
rect 3808 1760 4330 1761
rect 3808 1240 3809 1760
rect 4329 1240 4330 1760
rect 3808 1239 4330 1240
rect 2959 812 3063 1188
rect 2110 760 2632 761
rect 2110 240 2111 760
rect 2631 240 2632 760
rect 2110 239 2632 240
rect 1261 -188 1365 188
rect 412 -240 934 -239
rect 412 -760 413 -240
rect 933 -760 934 -240
rect 412 -761 934 -760
rect -437 -1188 -333 -812
rect -1286 -1240 -764 -1239
rect -1286 -1760 -1285 -1240
rect -765 -1760 -764 -1240
rect -1286 -1761 -764 -1760
rect -2135 -2000 -2031 -1812
rect -1077 -2000 -973 -1761
rect -437 -1812 -417 -1188
rect -353 -1812 -333 -1188
rect 621 -1239 725 -761
rect 1261 -812 1281 -188
rect 1345 -812 1365 -188
rect 2319 -239 2423 239
rect 2959 188 2979 812
rect 3043 188 3063 812
rect 4017 761 4121 1239
rect 4657 1188 4677 1812
rect 4741 1188 4761 1812
rect 5715 1761 5819 2000
rect 6355 1812 6459 2000
rect 5506 1760 6028 1761
rect 5506 1240 5507 1760
rect 6027 1240 6028 1760
rect 5506 1239 6028 1240
rect 4657 812 4761 1188
rect 3808 760 4330 761
rect 3808 240 3809 760
rect 4329 240 4330 760
rect 3808 239 4330 240
rect 2959 -188 3063 188
rect 2110 -240 2632 -239
rect 2110 -760 2111 -240
rect 2631 -760 2632 -240
rect 2110 -761 2632 -760
rect 1261 -1188 1365 -812
rect 412 -1240 934 -1239
rect 412 -1760 413 -1240
rect 933 -1760 934 -1240
rect 412 -1761 934 -1760
rect -437 -2000 -333 -1812
rect 621 -2000 725 -1761
rect 1261 -1812 1281 -1188
rect 1345 -1812 1365 -1188
rect 2319 -1239 2423 -761
rect 2959 -812 2979 -188
rect 3043 -812 3063 -188
rect 4017 -239 4121 239
rect 4657 188 4677 812
rect 4741 188 4761 812
rect 5715 761 5819 1239
rect 6355 1188 6375 1812
rect 6439 1188 6459 1812
rect 7413 1761 7517 2000
rect 8053 1812 8157 2000
rect 7204 1760 7726 1761
rect 7204 1240 7205 1760
rect 7725 1240 7726 1760
rect 7204 1239 7726 1240
rect 6355 812 6459 1188
rect 5506 760 6028 761
rect 5506 240 5507 760
rect 6027 240 6028 760
rect 5506 239 6028 240
rect 4657 -188 4761 188
rect 3808 -240 4330 -239
rect 3808 -760 3809 -240
rect 4329 -760 4330 -240
rect 3808 -761 4330 -760
rect 2959 -1188 3063 -812
rect 2110 -1240 2632 -1239
rect 2110 -1760 2111 -1240
rect 2631 -1760 2632 -1240
rect 2110 -1761 2632 -1760
rect 1261 -2000 1365 -1812
rect 2319 -2000 2423 -1761
rect 2959 -1812 2979 -1188
rect 3043 -1812 3063 -1188
rect 4017 -1239 4121 -761
rect 4657 -812 4677 -188
rect 4741 -812 4761 -188
rect 5715 -239 5819 239
rect 6355 188 6375 812
rect 6439 188 6459 812
rect 7413 761 7517 1239
rect 8053 1188 8073 1812
rect 8137 1188 8157 1812
rect 9111 1761 9215 2000
rect 9751 1812 9855 2000
rect 8902 1760 9424 1761
rect 8902 1240 8903 1760
rect 9423 1240 9424 1760
rect 8902 1239 9424 1240
rect 8053 812 8157 1188
rect 7204 760 7726 761
rect 7204 240 7205 760
rect 7725 240 7726 760
rect 7204 239 7726 240
rect 6355 -188 6459 188
rect 5506 -240 6028 -239
rect 5506 -760 5507 -240
rect 6027 -760 6028 -240
rect 5506 -761 6028 -760
rect 4657 -1188 4761 -812
rect 3808 -1240 4330 -1239
rect 3808 -1760 3809 -1240
rect 4329 -1760 4330 -1240
rect 3808 -1761 4330 -1760
rect 2959 -2000 3063 -1812
rect 4017 -2000 4121 -1761
rect 4657 -1812 4677 -1188
rect 4741 -1812 4761 -1188
rect 5715 -1239 5819 -761
rect 6355 -812 6375 -188
rect 6439 -812 6459 -188
rect 7413 -239 7517 239
rect 8053 188 8073 812
rect 8137 188 8157 812
rect 9111 761 9215 1239
rect 9751 1188 9771 1812
rect 9835 1188 9855 1812
rect 10809 1761 10913 2000
rect 11449 1812 11553 2000
rect 10600 1760 11122 1761
rect 10600 1240 10601 1760
rect 11121 1240 11122 1760
rect 10600 1239 11122 1240
rect 9751 812 9855 1188
rect 8902 760 9424 761
rect 8902 240 8903 760
rect 9423 240 9424 760
rect 8902 239 9424 240
rect 8053 -188 8157 188
rect 7204 -240 7726 -239
rect 7204 -760 7205 -240
rect 7725 -760 7726 -240
rect 7204 -761 7726 -760
rect 6355 -1188 6459 -812
rect 5506 -1240 6028 -1239
rect 5506 -1760 5507 -1240
rect 6027 -1760 6028 -1240
rect 5506 -1761 6028 -1760
rect 4657 -2000 4761 -1812
rect 5715 -2000 5819 -1761
rect 6355 -1812 6375 -1188
rect 6439 -1812 6459 -1188
rect 7413 -1239 7517 -761
rect 8053 -812 8073 -188
rect 8137 -812 8157 -188
rect 9111 -239 9215 239
rect 9751 188 9771 812
rect 9835 188 9855 812
rect 10809 761 10913 1239
rect 11449 1188 11469 1812
rect 11533 1188 11553 1812
rect 11449 812 11553 1188
rect 10600 760 11122 761
rect 10600 240 10601 760
rect 11121 240 11122 760
rect 10600 239 11122 240
rect 9751 -188 9855 188
rect 8902 -240 9424 -239
rect 8902 -760 8903 -240
rect 9423 -760 9424 -240
rect 8902 -761 9424 -760
rect 8053 -1188 8157 -812
rect 7204 -1240 7726 -1239
rect 7204 -1760 7205 -1240
rect 7725 -1760 7726 -1240
rect 7204 -1761 7726 -1760
rect 6355 -2000 6459 -1812
rect 7413 -2000 7517 -1761
rect 8053 -1812 8073 -1188
rect 8137 -1812 8157 -1188
rect 9111 -1239 9215 -761
rect 9751 -812 9771 -188
rect 9835 -812 9855 -188
rect 10809 -239 10913 239
rect 11449 188 11469 812
rect 11533 188 11553 812
rect 11449 -188 11553 188
rect 10600 -240 11122 -239
rect 10600 -760 10601 -240
rect 11121 -760 11122 -240
rect 10600 -761 11122 -760
rect 9751 -1188 9855 -812
rect 8902 -1240 9424 -1239
rect 8902 -1760 8903 -1240
rect 9423 -1760 9424 -1240
rect 8902 -1761 9424 -1760
rect 8053 -2000 8157 -1812
rect 9111 -2000 9215 -1761
rect 9751 -1812 9771 -1188
rect 9835 -1812 9855 -1188
rect 10809 -1239 10913 -761
rect 11449 -812 11469 -188
rect 11533 -812 11553 -188
rect 11449 -1188 11553 -812
rect 10600 -1240 11122 -1239
rect 10600 -1760 10601 -1240
rect 11121 -1760 11122 -1240
rect 10600 -1761 11122 -1760
rect 9751 -2000 9855 -1812
rect 10809 -2000 10913 -1761
rect 11449 -1812 11469 -1188
rect 11533 -1812 11553 -1188
rect 11449 -2000 11553 -1812
<< labels >>
rlabel via3 -10573 -1500 -10573 -1500 0 C2_0
port 1 nsew
rlabel mimcapcontact -11213 -1500 -11213 -1500 0 C1_0
port 2 nsew
rlabel via3 -8875 -1500 -8875 -1500 0 C2_1
port 3 nsew
rlabel mimcapcontact -9515 -1500 -9515 -1500 0 C1_1
port 4 nsew
rlabel via3 -7177 -1500 -7177 -1500 0 C2_2
port 5 nsew
rlabel mimcapcontact -7817 -1500 -7817 -1500 0 C1_2
port 6 nsew
rlabel via3 -5479 -1500 -5479 -1500 0 C2_3
port 7 nsew
rlabel mimcapcontact -6119 -1500 -6119 -1500 0 C1_3
port 8 nsew
rlabel via3 -3781 -1500 -3781 -1500 0 C2_4
port 9 nsew
rlabel mimcapcontact -4421 -1500 -4421 -1500 0 C1_4
port 10 nsew
rlabel via3 -2083 -1500 -2083 -1500 0 C2_5
port 11 nsew
rlabel mimcapcontact -2723 -1500 -2723 -1500 0 C1_5
port 12 nsew
rlabel via3 -385 -1500 -385 -1500 0 C2_6
port 13 nsew
rlabel mimcapcontact -1025 -1500 -1025 -1500 0 C1_6
port 14 nsew
rlabel via3 1313 -1500 1313 -1500 0 C2_7
port 15 nsew
rlabel mimcapcontact 673 -1500 673 -1500 0 C1_7
port 16 nsew
rlabel via3 3011 -1500 3011 -1500 0 C2_8
port 17 nsew
rlabel mimcapcontact 2371 -1500 2371 -1500 0 C1_8
port 18 nsew
rlabel via3 4709 -1500 4709 -1500 0 C2_9
port 19 nsew
rlabel mimcapcontact 4069 -1500 4069 -1500 0 C1_9
port 20 nsew
rlabel via3 6407 -1500 6407 -1500 0 C2_10
port 21 nsew
rlabel mimcapcontact 5767 -1500 5767 -1500 0 C1_10
port 22 nsew
rlabel via3 8105 -1500 8105 -1500 0 C2_11
port 23 nsew
rlabel mimcapcontact 7465 -1500 7465 -1500 0 C1_11
port 24 nsew
rlabel via3 9803 -1500 9803 -1500 0 C2_12
port 25 nsew
rlabel mimcapcontact 9163 -1500 9163 -1500 0 C1_12
port 26 nsew
rlabel via3 11501 -1500 11501 -1500 0 C2_13
port 27 nsew
rlabel mimcapcontact 10861 -1500 10861 -1500 0 C1_13
port 28 nsew
<< properties >>
string FIXED_BBOX 10521 1160 11201 1840
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 3.00 l 3.00 val 20.28 carea 2.00 cperi 0.19 class capacitor nx 14 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100 stack 1 doports 1
<< end >>
