magic
tech sky130A
magscale 1 2
timestamp 1762781875
<< metal1 >>
rect 27655 42880 47420 42890
rect 27655 42780 27665 42880
rect 27810 42780 47420 42880
rect 27655 42770 47420 42780
rect 27105 42225 46770 42235
rect 27105 42125 27115 42225
rect 27260 42125 46770 42225
rect 27105 42115 46770 42125
rect 26555 41570 46120 41580
rect 26555 41470 26565 41570
rect 26710 41470 46120 41570
rect 26555 41460 46120 41470
rect 26000 40920 45470 40930
rect 26000 40820 26010 40920
rect 26155 40820 45470 40920
rect 26000 40810 45470 40820
rect 45350 32335 45470 40810
rect 45350 32215 45855 32335
rect 7880 30260 14785 30665
rect 7880 1515 8285 30260
rect 45735 28840 45855 32215
rect 46000 30795 46120 41460
rect 46650 33410 46770 42115
rect 47300 34060 47420 42770
rect 47300 33940 55275 34060
rect 46650 33290 54680 33410
rect 45735 28740 45745 28840
rect 45845 28740 45855 28840
rect 45735 28730 45855 28740
rect 46000 27950 46120 27960
rect 46000 27850 46010 27950
rect 46110 27850 46120 27950
rect 46000 26620 46120 27850
rect 9585 25215 14785 25620
rect 9585 2555 9990 25215
rect 54560 22935 54680 33290
rect 45735 22815 54680 22935
rect 11290 22030 16235 22040
rect 11290 20865 11300 22030
rect 11930 20865 16235 22030
rect 11290 20855 16235 20865
rect 11290 19560 14785 19965
rect 11290 3625 11695 19560
rect 45735 18140 45855 22815
rect 55155 22340 55275 33940
rect 46000 22220 55275 22340
rect 46000 20095 46120 22220
rect 45735 18040 45745 18140
rect 45845 18040 45855 18140
rect 45735 18030 45855 18040
rect 46000 17250 46120 17260
rect 46000 17150 46010 17250
rect 46110 17150 46120 17250
rect 46000 15925 46120 17150
rect 12995 14515 14785 14920
rect 12995 4680 13400 14515
rect 12995 4670 26680 4680
rect 12995 4285 26285 4670
rect 26670 4285 26680 4670
rect 12995 4275 26680 4285
rect 11290 3615 22815 3625
rect 11290 3230 22420 3615
rect 22805 3230 22815 3615
rect 11290 3220 22815 3230
rect 9585 2545 18950 2555
rect 9585 2160 18555 2545
rect 18940 2160 18950 2545
rect 9585 2150 18950 2160
rect 7880 1505 15085 1515
rect 7880 1140 14690 1505
rect 15075 1140 15085 1505
rect 7880 1130 15085 1140
<< via1 >>
rect 27665 42780 27810 42880
rect 27115 42125 27260 42225
rect 26565 41470 26710 41570
rect 26010 40820 26155 40920
rect 45745 28740 45845 28840
rect 46010 27850 46110 27950
rect 11300 20865 11930 22030
rect 45745 18040 45845 18140
rect 46010 17150 46110 17250
rect 26285 4285 26670 4670
rect 22420 3230 22805 3615
rect 18555 2160 18940 2545
rect 14690 1140 15075 1505
<< metal2 >>
rect 11290 43420 25520 43430
rect 11290 43030 25300 43420
rect 25510 43030 25520 43420
rect 11290 43020 25520 43030
rect 11290 27450 11695 43020
rect 27655 42880 27820 42890
rect 27655 42780 27665 42880
rect 27810 42780 27820 42880
rect 27655 42770 27820 42780
rect 27105 42225 27270 42235
rect 27105 42125 27115 42225
rect 27260 42125 27270 42225
rect 27105 42115 27270 42125
rect 26555 41570 26720 41580
rect 26555 41470 26565 41570
rect 26710 41470 26720 41570
rect 26555 41460 26720 41470
rect 26000 40920 26165 40930
rect 26000 40820 26010 40920
rect 26155 40820 26165 40920
rect 26000 40810 26165 40820
rect 45735 28840 45855 28850
rect 45735 28740 45745 28840
rect 45845 28740 45855 28840
rect 45735 27960 45855 28740
rect 45735 27950 46120 27960
rect 45735 27850 46010 27950
rect 46110 27850 46120 27950
rect 45735 27840 46120 27850
rect 11290 27200 14535 27450
rect 11290 22030 16235 22040
rect 11290 20865 11300 22030
rect 11930 20865 16235 22030
rect 11290 20855 16235 20865
rect 45735 18140 45855 18150
rect 45735 18040 45745 18140
rect 45845 18040 45855 18140
rect 45735 17260 45855 18040
rect 45735 17250 46120 17260
rect 45735 17150 46010 17250
rect 46110 17150 46120 17250
rect 45735 17140 46120 17150
rect 26275 4670 26680 4680
rect 26275 4285 26285 4670
rect 26670 4285 26680 4670
rect 26275 4275 26680 4285
rect 22410 3615 22815 3625
rect 22410 3230 22420 3615
rect 22805 3230 22815 3615
rect 22410 3220 22815 3230
rect 18545 2545 18950 2555
rect 18545 2160 18555 2545
rect 18940 2160 18950 2545
rect 18545 2150 18950 2160
rect 14680 1505 15085 1515
rect 14680 1140 14690 1505
rect 15075 1140 15085 1505
rect 14680 1130 15085 1140
<< via2 >>
rect 25300 43030 25510 43420
rect 27665 42780 27810 42880
rect 27115 42125 27260 42225
rect 26565 41470 26710 41570
rect 26010 40820 26155 40920
rect 11300 20865 11930 22030
rect 26285 4285 26670 4670
rect 22420 3230 22805 3615
rect 18555 2160 18940 2545
rect 14690 1140 15075 1505
<< metal3 >>
rect 25290 43420 25520 43430
rect 25290 43030 25300 43420
rect 25510 43030 25520 43420
rect 25290 43020 25520 43030
rect 27655 42880 27820 42890
rect 27655 42780 27665 42880
rect 27810 42780 27820 42880
rect 27655 42770 27820 42780
rect 27105 42225 27270 42235
rect 27105 42125 27115 42225
rect 27260 42125 27270 42225
rect 27105 42115 27270 42125
rect 26555 41570 26720 41580
rect 26555 41470 26565 41570
rect 26710 41470 26720 41570
rect 26555 41460 26720 41470
rect 26000 40920 26165 40930
rect 26000 40820 26010 40920
rect 26155 40820 26165 40920
rect 26000 40810 26165 40820
rect 200 25865 13000 25875
rect 200 24700 210 25865
rect 590 24700 13000 25865
rect 200 24690 13000 24700
rect 800 22030 11940 22040
rect 800 20865 810 22030
rect 1190 20865 11300 22030
rect 11930 20865 11940 22030
rect 800 20855 11940 20865
rect 26275 4670 26680 4680
rect 26275 4285 26285 4670
rect 26670 4285 26680 4670
rect 26275 4275 26680 4285
rect 22410 3615 22815 3625
rect 22410 3230 22420 3615
rect 22805 3230 22815 3615
rect 22410 3220 22815 3230
rect 18545 2545 18950 2555
rect 18545 2160 18555 2545
rect 18940 2160 18950 2545
rect 18545 2150 18950 2160
rect 54420 1740 55030 14280
rect 30360 1730 55030 1740
rect 14680 1505 15085 1515
rect 14680 1140 14690 1505
rect 15075 1140 15085 1505
rect 14680 1130 15085 1140
rect 30360 1140 30370 1730
rect 30945 1140 55030 1730
rect 30360 1130 55030 1140
<< via3 >>
rect 25300 43030 25510 43420
rect 27665 42780 27810 42880
rect 27115 42125 27260 42225
rect 26565 41470 26710 41570
rect 26010 40820 26155 40920
rect 210 24700 590 25865
rect 810 20865 1190 22030
rect 26285 4285 26670 4670
rect 22420 3230 22805 3615
rect 18555 2160 18940 2545
rect 14690 1140 15075 1505
rect 30370 1140 30945 1730
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 44952 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 45060 25514 45152
rect 26006 45060 26066 45152
rect 26558 45060 26618 45152
rect 27110 45060 27170 45152
rect 27662 45060 27722 45152
rect 200 25865 600 44152
rect 200 24700 210 25865
rect 590 24700 600 25865
rect 200 1000 600 24700
rect 800 22030 1200 44152
rect 25450 43430 25520 45060
rect 25290 43420 25520 43430
rect 25290 43030 25300 43420
rect 25510 43030 25520 43420
rect 25290 43020 25520 43030
rect 26000 40930 26070 45060
rect 26555 41580 26625 45060
rect 27105 42235 27175 45060
rect 27655 42890 27725 45060
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 27655 42880 27820 42890
rect 27655 42780 27665 42880
rect 27810 42780 27820 42880
rect 27655 42770 27820 42780
rect 27105 42225 27270 42235
rect 27105 42125 27115 42225
rect 27260 42125 27270 42225
rect 27105 42115 27270 42125
rect 26555 41570 26720 41580
rect 26555 41470 26565 41570
rect 26710 41470 26720 41570
rect 26555 41460 26720 41470
rect 26000 40920 26165 40930
rect 26000 40820 26010 40920
rect 26155 40820 26165 40920
rect 26000 40810 26165 40820
rect 800 20865 810 22030
rect 1190 20865 1200 22030
rect 800 1000 1200 20865
rect 26275 4670 26680 4680
rect 26275 4285 26285 4670
rect 26670 4285 26680 4670
rect 22410 3615 22815 3625
rect 22410 3230 22420 3615
rect 22805 3230 22815 3615
rect 18545 2545 18950 2555
rect 18545 2160 18555 2545
rect 18940 2160 18950 2545
rect 14680 1505 15085 1515
rect 14680 1140 14690 1505
rect 15075 1140 15085 1505
rect 14680 1130 15085 1140
rect 18545 1130 18950 2160
rect 22410 1130 22815 3230
rect 26275 1130 26680 4285
rect 14905 200 15085 1130
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 1130
rect 22630 200 22815 1130
rect 26495 200 26680 1130
rect 30360 1730 30955 1740
rect 30360 1140 30370 1730
rect 30945 1140 30955 1730
rect 30360 1130 30955 1140
rect 30360 200 30545 1130
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30362 0 30542 200
<< comment >>
rect 63600 44600 66800 45000
rect 66400 400 66800 44600
rect 63600 0 66800 400
use iq_modulator  iq_modulator_0
timestamp 1762715922
transform 1 0 18600 0 1 20200
box -5600 -15200 36430 20020
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 66976 45152
<< end >>
