magic
tech sky130A
magscale 1 2
timestamp 1762641840
<< locali >>
rect -130 4680 2270 4695
rect -130 4555 -115 4680
rect 2255 4555 2270 4680
rect -130 4395 325 4555
rect 1810 4395 2270 4555
rect -130 4260 2270 4395
rect -130 4065 25 4260
rect -130 2290 -100 4065
rect -60 2290 25 4065
rect -130 2155 25 2290
rect 2115 4065 2270 4260
rect 2115 2290 2195 4065
rect 2235 2290 2270 4065
rect 2115 2155 2270 2290
rect -130 2130 2270 2155
rect -130 2095 25 2130
rect 2115 2095 2270 2130
rect -130 1925 2270 1985
rect -130 1800 25 1925
rect -130 1220 -100 1800
rect -60 1220 25 1800
rect -130 1070 25 1220
rect 2115 1800 2270 1925
rect 2115 1220 2195 1800
rect 2235 1220 2270 1800
rect 2115 1070 2270 1220
rect -130 905 2270 1070
rect -130 745 325 905
rect 1810 745 2270 905
rect -130 620 -115 745
rect 2255 620 2270 745
rect -130 605 2270 620
<< viali >>
rect -115 4555 2255 4680
rect 325 4395 1810 4555
rect -100 2290 -60 4065
rect 2195 2290 2235 4065
rect -100 1220 -60 1800
rect 2195 1220 2235 1800
rect 325 745 1810 905
rect -115 620 2255 745
<< metal1 >>
rect -130 4680 2270 4695
rect -130 4555 -115 4680
rect 2255 4555 2270 4680
rect -130 4540 325 4555
rect -130 4080 20 4540
rect 70 4435 240 4450
rect 70 4315 85 4435
rect 225 4315 240 4435
rect 310 4395 325 4540
rect 1810 4540 2270 4555
rect 1810 4395 1825 4540
rect 310 4380 1825 4395
rect 1895 4435 2065 4450
rect 70 4130 240 4315
rect 1895 4315 1910 4435
rect 2050 4315 2065 4435
rect 290 4135 1845 4295
rect 290 4080 380 4135
rect -130 4065 235 4080
rect -130 2290 -100 4065
rect -60 2290 85 4065
rect 225 2290 235 4065
rect -130 2275 235 2290
rect 270 2275 380 4080
rect 475 4070 635 4080
rect 475 2285 485 4070
rect 625 2285 635 4070
rect 475 2275 635 2285
rect 730 2275 890 4135
rect 990 4070 1150 4080
rect 990 2285 1000 4070
rect 1140 2285 1150 4070
rect 990 2275 1150 2285
rect 1250 2275 1410 4135
rect 1760 4080 1845 4135
rect 1895 4130 2065 4315
rect 2115 4080 2270 4540
rect 1505 4070 1665 4080
rect 1505 2285 1515 4070
rect 1655 2285 1665 4070
rect 1505 2275 1665 2285
rect 1760 2275 1920 4080
rect 2085 4065 2270 4080
rect 2085 2290 2195 4065
rect 2235 2290 2270 4065
rect 2085 2275 2270 2290
rect 730 2230 890 2235
rect 330 2195 1810 2230
rect -165 1885 1810 2195
rect 330 1850 1810 1885
rect 730 1845 890 1850
rect -130 1810 60 1815
rect -130 1800 55 1810
rect -130 1220 -100 1800
rect -60 1220 55 1800
rect -130 1205 55 1220
rect 215 1210 375 1810
rect 475 1800 635 1810
rect 475 1220 485 1800
rect 625 1220 635 1800
rect 475 1210 635 1220
rect -130 760 20 1205
rect 70 985 240 1170
rect 290 1155 375 1210
rect 730 1155 890 1810
rect 990 1800 1150 1810
rect 990 1220 1000 1800
rect 1140 1220 1150 1800
rect 990 1210 1150 1220
rect 1245 1155 1405 1810
rect 1505 1800 1665 1810
rect 1505 1220 1515 1800
rect 1655 1220 1665 1800
rect 1505 1210 1665 1220
rect 1760 1210 1920 1810
rect 2085 1800 2270 1815
rect 2085 1220 2195 1800
rect 2235 1220 2270 1800
rect 2085 1210 2270 1220
rect 1760 1155 1845 1210
rect 290 995 1845 1155
rect 70 865 85 985
rect 225 865 240 985
rect 1895 985 2065 1170
rect 70 850 240 865
rect 310 905 1825 920
rect 310 760 325 905
rect -130 745 325 760
rect 1810 760 1825 905
rect 1895 865 1910 985
rect 2050 865 2065 985
rect 1895 850 2065 865
rect 2115 760 2270 1210
rect 1810 745 2270 760
rect -130 620 -115 745
rect 2255 620 2270 745
rect -130 605 2270 620
<< via1 >>
rect 85 4315 225 4435
rect 1910 4315 2050 4435
rect 85 2290 225 4065
rect 485 2285 625 4070
rect 1000 2285 1140 4070
rect 1515 2285 1655 4070
rect 485 1220 625 1800
rect 1000 1220 1140 1800
rect 1515 1220 1655 1800
rect 85 865 225 985
rect 1910 865 2050 985
<< metal2 >>
rect -165 4435 2065 4450
rect -165 4315 85 4435
rect 225 4315 1910 4435
rect 2050 4315 2065 4435
rect -165 4300 2065 4315
rect 70 4065 240 4080
rect 70 2290 85 4065
rect 225 2290 240 4065
rect 70 1000 240 2290
rect 475 4070 635 4080
rect 475 2285 485 4070
rect 625 2285 635 4070
rect 475 2240 635 2285
rect 990 4070 1150 4080
rect 990 2285 1000 4070
rect 1140 2285 1150 4070
rect 990 2240 1150 2285
rect 1505 4070 1665 4080
rect 1505 2285 1515 4070
rect 1655 2285 1665 4070
rect 1505 2240 1665 2285
rect 475 1840 2305 2240
rect 475 1800 635 1840
rect 475 1220 485 1800
rect 625 1220 635 1800
rect 475 1210 635 1220
rect 990 1800 1150 1840
rect 990 1220 1000 1800
rect 1140 1220 1150 1800
rect 990 1210 1150 1220
rect 1505 1800 1665 1840
rect 1505 1220 1515 1800
rect 1655 1220 1665 1800
rect 1505 1210 1665 1220
rect 70 985 2065 1000
rect 70 865 85 985
rect 225 865 1910 985
rect 2050 865 2065 985
rect 70 850 2065 865
use sky130_fd_pr__nfet_01v8_lvt_WHJEU4  sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0
timestamp 1762641840
transform 1 0 1069 0 1 1510
box -1199 -510 1199 510
use sky130_fd_pr__pfet_01v8_lvt_P4QH36  sky130_fd_pr__pfet_01v8_lvt_P4QH36_0
timestamp 1762641840
transform 1 0 1069 0 1 3179
box -1199 -1119 1199 1119
<< labels >>
flabel metal2 -155 4370 -155 4370 0 FreeSans 320 0 0 0 di_en
port 8 nsew
flabel viali 1040 670 1040 670 0 FreeSans 400 0 0 0 VSS
port 10 nsew
flabel metal1 -155 2040 -155 2040 0 FreeSans 320 0 0 0 vin
port 12 nsew
flabel metal2 2265 2035 2265 2035 0 FreeSans 320 0 0 0 vout
port 13 nsew
flabel viali 965 4610 965 4610 0 FreeSans 400 0 0 0 VDD
port 11 nsew
<< end >>
