magic
tech sky130A
magscale 1 2
timestamp 1762090404
<< metal1 >>
rect 8430 6945 8650 7350
rect -2685 6680 2385 6805
rect -2680 2970 -2345 6680
rect -2105 6145 2510 6550
rect 5275 6145 5500 6550
rect 25435 6530 25715 6550
rect 18870 6500 18960 6505
rect 25435 6165 25470 6530
rect 25695 6165 25715 6530
rect 25435 6145 25715 6165
rect -2155 5715 -1930 5865
rect -2105 3155 -2055 3265
rect -2680 2390 -1970 2970
rect -2225 1775 -1905 1925
rect -2110 1100 2510 1505
rect 5280 1100 5495 1505
rect 25450 1485 25715 1505
rect 25450 1120 25470 1485
rect 25695 1120 25715 1485
rect 25450 1100 25715 1120
rect 8430 300 8650 705
<< via1 >>
rect 18870 6185 18960 6500
rect 25470 6165 25695 6530
rect 2260 1790 2370 1910
rect 18870 1145 18960 1460
rect 25470 1120 25695 1485
rect 2295 855 2370 950
<< metal2 >>
rect 25450 6530 25715 6550
rect 18855 6500 18975 6515
rect 18855 6185 18870 6500
rect 18960 6185 18975 6500
rect 18855 6170 18975 6185
rect 25450 6165 25470 6530
rect 25695 6165 25715 6530
rect 25450 6145 25715 6165
rect -135 5470 60 5620
rect 2245 1910 2385 1925
rect 2245 1790 2260 1910
rect 2370 1790 2385 1910
rect 2245 950 2385 1790
rect 25450 1485 25715 1505
rect 18855 1460 18975 1475
rect 18855 1145 18870 1460
rect 18960 1145 18975 1460
rect 18855 1130 18975 1145
rect 25450 1120 25470 1485
rect 25695 1120 25715 1485
rect 25450 1100 25715 1120
rect 2245 855 2295 950
rect 2370 855 2385 950
rect 2245 840 2385 855
<< via2 >>
rect 18870 6185 18960 6500
rect 25470 6165 25695 6530
rect 18870 1145 18960 1460
rect 25470 1120 25695 1485
<< metal3 >>
rect 25450 6530 28500 6550
rect 7375 6500 18975 6515
rect 7375 6185 18870 6500
rect 18960 6185 18975 6500
rect 7375 6170 18975 6185
rect 7375 5960 7540 6170
rect 25450 6165 25470 6530
rect 25695 6165 28500 6530
rect 25450 5965 28500 6165
rect -2105 5615 7540 5960
rect 10010 5615 28500 5965
rect -2105 1685 10205 2020
rect 12675 1685 28500 2020
rect 10035 1475 10205 1685
rect 25450 1485 28500 1685
rect 10035 1460 18975 1475
rect 10035 1145 18870 1460
rect 18960 1145 18975 1460
rect 10035 1130 18975 1145
rect 25450 1120 25470 1485
rect 25695 1120 28500 1485
rect 25450 1100 28500 1120
use ota_core_hybrid_bm  ota_core_hybrid_bm_0 ota_core
timestamp 1761868878
transform 1 0 3061 0 1 94
box -5165 1680 25175 5770
use resistors  resistors_0 resistors
timestamp 1761785752
transform 1 0 2310 0 1 -1385
box -65 1425 23150 8995
<< labels >>
flabel metal1 -1914 6358 -1914 6358 0 FreeSans 1200 0 0 0 vinp
port 3 nsew
flabel metal1 -1916 1306 -1916 1306 0 FreeSans 1200 0 0 0 vinn
port 5 nsew
flabel metal1 -2135 5790 -2135 5790 0 FreeSans 800 0 0 0 VDD
port 10 nsew
flabel metal1 -2175 1850 -2175 1850 0 FreeSans 800 0 0 0 VSS
port 11 nsew
flabel metal1 5385 6360 5385 6360 0 FreeSans 400 0 0 0 vC1p
port 29 nsew
flabel metal1 5380 1305 5380 1305 0 FreeSans 400 0 0 0 vC1n
port 31 nsew
flabel metal1 8530 590 8530 590 0 FreeSans 400 0 0 0 vC2n
port 33 nsew
flabel metal1 8540 7150 8540 7150 0 FreeSans 400 0 0 0 vC2p
port 35 nsew
flabel metal1 -2080 3205 -2080 3205 0 FreeSans 400 0 0 0 di_filter_ota_en
port 37 nsew
flabel metal3 28190 6150 28190 6150 0 FreeSans 1200 0 0 0 voutn
port 46 nsew
flabel metal3 28220 1505 28220 1505 0 FreeSans 1200 0 0 0 voutp
port 48 nsew
<< end >>
