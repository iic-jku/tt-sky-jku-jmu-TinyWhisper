magic
tech sky130A
magscale 1 2
timestamp 1762800247
<< locali >>
rect 7150 30250 15060 31970
rect 7150 30115 15055 30250
rect 7145 23210 15060 25760
rect 7145 20870 11305 23210
rect 11925 20870 15060 23210
rect 7145 19415 15060 20870
rect 7150 13190 15055 15060
<< viali >>
rect 11305 20870 11925 23210
rect 15070 21940 16220 22245
<< metal1 >>
rect 800 40760 1605 43055
rect 27655 42880 47420 42890
rect 3500 42805 6505 42815
rect 3500 42750 3510 42805
rect 6495 42750 6505 42805
rect 27655 42780 27665 42880
rect 27810 42780 47420 42880
rect 27655 42770 47420 42780
rect 3500 42740 6505 42750
rect 27105 42225 46770 42235
rect 27105 42125 27115 42225
rect 27260 42125 46770 42225
rect 27105 42115 46770 42125
rect 26555 41570 46120 41580
rect 26555 41470 26565 41570
rect 26710 41470 46120 41570
rect 26555 41460 46120 41470
rect 26000 40920 45470 40930
rect 26000 40820 26010 40920
rect 26155 40820 45470 40920
rect 26000 40810 45470 40820
rect 800 40720 7040 40760
rect 800 39980 840 40720
rect 1160 39980 7040 40720
rect 800 39940 7040 39980
rect 800 35620 1605 39940
rect 2995 37550 6995 37705
rect 800 35580 7020 35620
rect 800 34840 840 35580
rect 1160 34840 7020 35580
rect 800 34800 7020 34840
rect 800 31600 1605 34800
rect 2995 32330 6995 32490
rect 45350 32335 45470 40810
rect 45350 32215 45855 32335
rect 800 31360 840 31600
rect 1160 31360 1605 31600
rect 800 30080 1605 31360
rect 7880 30260 14785 30665
rect 800 29260 7040 30080
rect 800 28800 1605 29260
rect 800 28060 840 28800
rect 1160 28060 1605 28800
rect 800 25160 1605 28060
rect 2995 27110 6995 27270
rect 800 24340 7020 25160
rect 800 23180 1605 24340
rect 800 20900 840 23180
rect 1160 20900 1605 23180
rect 2995 21895 6995 22050
rect 800 19820 1605 20900
rect 800 19000 7020 19820
rect 800 14620 1605 19000
rect 2995 16675 6995 16835
rect 800 13820 7020 14620
rect 800 13580 840 13820
rect 1160 13800 7020 13820
rect 1160 13580 1605 13800
rect 800 9360 1605 13580
rect 2995 11460 6995 11615
rect 800 9320 7020 9360
rect 800 8580 840 9320
rect 1160 8580 7020 9320
rect 800 8540 7020 8580
rect 800 4160 1605 8540
rect 2995 6240 6995 6400
rect 800 4120 7020 4160
rect 800 3380 840 4120
rect 1160 3380 7020 4120
rect 800 3340 7020 3380
rect 800 1035 1605 3340
rect 7880 1515 8285 30260
rect 45735 28840 45855 32215
rect 46000 30795 46120 41460
rect 46650 33410 46770 42115
rect 47300 34060 47420 42770
rect 47300 33940 55275 34060
rect 46650 33290 54680 33410
rect 45735 28740 45745 28840
rect 45845 28740 45855 28840
rect 45735 28730 45855 28740
rect 46000 27950 46120 27960
rect 46000 27850 46010 27950
rect 46110 27850 46120 27950
rect 46000 26620 46120 27850
rect 9585 25215 14785 25620
rect 9585 2555 9990 25215
rect 15055 23225 16235 24570
rect 11290 23215 16235 23225
rect 11290 20865 11300 23215
rect 11930 22245 16235 23215
rect 54560 22935 54680 33290
rect 11930 21940 15070 22245
rect 16220 21940 16235 22245
rect 11930 20865 16235 21940
rect 11290 20855 16235 20865
rect 15055 20610 16235 20855
rect 45735 22815 54680 22935
rect 11290 19560 14785 19965
rect 11290 3625 11695 19560
rect 45735 18140 45855 22815
rect 55155 22340 55275 33940
rect 46000 22220 55275 22340
rect 46000 20095 46120 22220
rect 45735 18040 45745 18140
rect 45845 18040 45855 18140
rect 45735 18030 45855 18040
rect 46000 17250 46120 17260
rect 46000 17150 46010 17250
rect 46110 17150 46120 17250
rect 46000 15925 46120 17150
rect 12995 14515 14785 14920
rect 12995 4680 13400 14515
rect 12995 4670 26680 4680
rect 12995 4285 26285 4670
rect 26670 4285 26680 4670
rect 12995 4275 26680 4285
rect 11290 3615 22815 3625
rect 11290 3230 22420 3615
rect 22805 3230 22815 3615
rect 11290 3220 22815 3230
rect 9585 2545 18950 2555
rect 9585 2160 18555 2545
rect 18940 2160 18950 2545
rect 9585 2150 18950 2160
rect 7880 1505 15085 1515
rect 3490 1195 6505 1205
rect 3490 1180 3500 1195
rect 2995 1140 3500 1180
rect 6495 1180 6505 1195
rect 6495 1140 6995 1180
rect 2995 1130 6995 1140
rect 7880 1140 14690 1505
rect 15075 1140 15085 1505
rect 7880 1130 15085 1140
<< via1 >>
rect 3510 42750 6495 42805
rect 27665 42780 27810 42880
rect 27115 42125 27260 42225
rect 26565 41470 26710 41570
rect 26010 40820 26155 40920
rect 840 39980 1160 40720
rect 840 34840 1160 35580
rect 840 31360 1160 31600
rect 840 28060 1160 28800
rect 840 20900 1160 23180
rect 840 13580 1160 13820
rect 840 8580 1160 9320
rect 840 3380 1160 4120
rect 45745 28740 45845 28840
rect 46010 27850 46110 27950
rect 11300 23210 11930 23215
rect 11300 20870 11305 23210
rect 11305 20870 11925 23210
rect 11925 20870 11930 23210
rect 11300 20865 11930 20870
rect 45745 18040 45845 18140
rect 46010 17150 46110 17250
rect 26285 4285 26670 4670
rect 22420 3230 22805 3615
rect 18555 2160 18940 2545
rect 3500 1140 6495 1195
rect 14690 1140 15075 1505
<< metal2 >>
rect 11290 43420 25520 43430
rect 11290 43030 25300 43420
rect 25510 43030 25520 43420
rect 11290 43020 25520 43030
rect 3500 42805 6505 42815
rect 3500 42750 3510 42805
rect 6495 42750 6505 42805
rect 800 40720 1200 40760
rect 800 39980 840 40720
rect 1160 39980 1200 40720
rect 800 39940 1200 39980
rect 800 35580 1200 35620
rect 800 34840 840 35580
rect 1160 34840 1200 35580
rect 800 34800 1200 34840
rect 800 31600 1200 31640
rect 800 31360 840 31600
rect 1160 31360 1200 31600
rect 800 31320 1200 31360
rect 3500 29970 6505 42750
rect 6495 29645 6505 29970
rect 800 28800 1200 28840
rect 800 28060 840 28800
rect 1160 28060 1200 28800
rect 800 28020 1200 28060
rect 3500 25865 6505 29645
rect 11290 27450 11695 43020
rect 27655 42880 27820 42890
rect 27655 42780 27665 42880
rect 27810 42780 27820 42880
rect 27655 42770 27820 42780
rect 27105 42225 27270 42235
rect 27105 42125 27115 42225
rect 27260 42125 27270 42225
rect 27105 42115 27270 42125
rect 26555 41570 26720 41580
rect 26555 41470 26565 41570
rect 26710 41470 26720 41570
rect 26555 41460 26720 41470
rect 26000 40920 26165 40930
rect 26000 40820 26010 40920
rect 26155 40820 26165 40920
rect 26000 40810 26165 40820
rect 45735 28840 45855 28850
rect 45735 28740 45745 28840
rect 45845 28740 45855 28840
rect 45735 27960 45855 28740
rect 45735 27950 46120 27960
rect 45735 27850 46010 27950
rect 46110 27850 46120 27950
rect 45735 27840 46120 27850
rect 11290 27200 14535 27450
rect 6495 24700 6505 25865
rect 800 23180 1200 23220
rect 800 20900 840 23180
rect 1160 20900 1200 23180
rect 800 20860 1200 20900
rect 3500 19270 6505 24700
rect 15055 23225 16235 24570
rect 11290 23215 16235 23225
rect 11290 20865 11300 23215
rect 11930 20865 16235 23215
rect 11290 20855 16235 20865
rect 15055 20610 16235 20855
rect 6495 18945 6505 19270
rect 800 13820 1200 13860
rect 800 13580 840 13820
rect 1160 13580 1200 13820
rect 800 13540 1200 13580
rect 800 9320 1200 9360
rect 800 8580 840 9320
rect 1160 8580 1200 9320
rect 800 8540 1200 8580
rect 800 4120 1200 4160
rect 800 3380 840 4120
rect 1160 3380 1200 4120
rect 800 3340 1200 3380
rect 3500 1205 6505 18945
rect 45735 18140 45855 18150
rect 45735 18040 45745 18140
rect 45845 18040 45855 18140
rect 45735 17260 45855 18040
rect 45735 17250 46120 17260
rect 45735 17150 46010 17250
rect 46110 17150 46120 17250
rect 45735 17140 46120 17150
rect 26275 4670 26680 4680
rect 26275 4285 26285 4670
rect 26670 4285 26680 4670
rect 26275 4275 26680 4285
rect 22410 3615 22815 3625
rect 22410 3230 22420 3615
rect 22805 3230 22815 3615
rect 22410 3220 22815 3230
rect 18545 2545 18950 2555
rect 18545 2160 18555 2545
rect 18940 2160 18950 2545
rect 18545 2150 18950 2160
rect 3490 1195 6505 1205
rect 3490 1140 3500 1195
rect 6495 1140 6505 1195
rect 3490 1130 6505 1140
rect 14680 1505 15085 1515
rect 14680 1140 14690 1505
rect 15075 1140 15085 1505
rect 14680 1130 15085 1140
<< via2 >>
rect 25300 43030 25510 43420
rect 840 39980 1160 40720
rect 840 34840 1160 35580
rect 840 31360 1160 31600
rect 3500 29645 6495 29970
rect 840 28060 1160 28800
rect 27665 42780 27810 42880
rect 27115 42125 27260 42225
rect 26565 41470 26710 41570
rect 26010 40820 26155 40920
rect 3500 24700 6495 25865
rect 840 20900 1160 23180
rect 11300 20865 11930 23215
rect 3500 18945 6495 19270
rect 840 13580 1160 13820
rect 840 8580 1160 9320
rect 840 3380 1160 4120
rect 26285 4285 26670 4670
rect 22420 3230 22805 3615
rect 18555 2160 18940 2545
rect 14690 1140 15075 1505
<< metal3 >>
rect 25290 43420 25520 43430
rect 25290 43030 25300 43420
rect 25510 43030 25520 43420
rect 25290 43020 25520 43030
rect 27655 42880 27820 42890
rect 27655 42780 27665 42880
rect 27810 42780 27820 42880
rect 27655 42770 27820 42780
rect 27105 42225 27270 42235
rect 27105 42125 27115 42225
rect 27260 42125 27270 42225
rect 27105 42115 27270 42125
rect 26555 41570 26720 41580
rect 26555 41470 26565 41570
rect 26710 41470 26720 41570
rect 26555 41460 26720 41470
rect 26000 40920 26165 40930
rect 26000 40820 26010 40920
rect 26155 40820 26165 40920
rect 26000 40810 26165 40820
rect 800 40720 1200 40760
rect 800 39980 840 40720
rect 1160 39980 1200 40720
rect 800 39940 1200 39980
rect 800 35580 1200 35620
rect 800 34840 840 35580
rect 1160 34840 1200 35580
rect 800 34800 1200 34840
rect 800 31635 15060 31645
rect 800 31320 810 31635
rect 1190 31320 15060 31635
rect 800 31310 15060 31320
rect 200 29970 13000 29980
rect 200 29645 210 29970
rect 590 29645 3500 29970
rect 6495 29645 13000 29970
rect 200 29635 13000 29645
rect 800 28800 1200 28840
rect 800 28060 840 28800
rect 1160 28060 1200 28800
rect 800 28020 1200 28060
rect 200 25865 13000 25875
rect 200 24700 210 25865
rect 590 24700 3500 25865
rect 6495 24700 13000 25865
rect 200 24690 13000 24700
rect 800 23215 11940 23225
rect 800 20865 810 23215
rect 1190 20865 11300 23215
rect 11930 20865 11940 23215
rect 800 20855 11940 20865
rect 200 19270 13005 19280
rect 200 18945 210 19270
rect 590 18945 3500 19270
rect 6495 18945 13005 19270
rect 200 18935 13005 18945
rect 800 13860 15060 13870
rect 800 13545 810 13860
rect 1190 13545 15060 13860
rect 800 13535 15060 13545
rect 800 9320 1200 9360
rect 800 8580 840 9320
rect 1160 8580 1200 9320
rect 800 8540 1200 8580
rect 26275 4670 26680 4680
rect 26275 4285 26285 4670
rect 26670 4285 26680 4670
rect 26275 4275 26680 4285
rect 800 4120 1200 4160
rect 800 3380 840 4120
rect 1160 3380 1200 4120
rect 800 3340 1200 3380
rect 22410 3615 22815 3625
rect 22410 3230 22420 3615
rect 22805 3230 22815 3615
rect 22410 3220 22815 3230
rect 18545 2545 18950 2555
rect 18545 2160 18555 2545
rect 18940 2160 18950 2545
rect 18545 2150 18950 2160
rect 54420 1740 55030 14280
rect 30360 1730 55030 1740
rect 14680 1505 15085 1515
rect 14680 1140 14690 1505
rect 15075 1140 15085 1505
rect 14680 1130 15085 1140
rect 30360 1140 30370 1730
rect 30945 1140 55030 1730
rect 30360 1130 55030 1140
<< via3 >>
rect 25300 43030 25510 43420
rect 27665 42780 27810 42880
rect 27115 42125 27260 42225
rect 26565 41470 26710 41570
rect 26010 40820 26155 40920
rect 840 39980 1160 40720
rect 840 34840 1160 35580
rect 52675 31715 53265 31955
rect 810 31600 1190 31635
rect 810 31360 840 31600
rect 840 31360 1160 31600
rect 1160 31360 1190 31600
rect 810 31320 1190 31360
rect 210 29645 590 29970
rect 840 28060 1160 28800
rect 51685 28075 52275 28315
rect 210 24700 590 25865
rect 810 23180 1190 23215
rect 810 20900 840 23180
rect 840 20900 1160 23180
rect 1160 20900 1190 23180
rect 810 20865 1190 20900
rect 210 18945 590 19270
rect 51685 17375 52275 17615
rect 52675 16845 53265 17085
rect 810 13820 1190 13860
rect 810 13580 840 13820
rect 840 13580 1160 13820
rect 1160 13580 1190 13820
rect 810 13545 1190 13580
rect 840 8580 1160 9320
rect 26285 4285 26670 4670
rect 840 3380 1160 4120
rect 22420 3230 22805 3615
rect 18555 2160 18940 2545
rect 14690 1140 15075 1505
rect 30370 1140 30945 1730
<< metal4 >>
rect 6134 45065 6194 45152
rect 6686 45065 6746 45152
rect 7238 45065 7298 45152
rect 7790 45065 7850 45152
rect 8342 45065 8402 45152
rect 8894 45065 8954 45152
rect 9446 45065 9506 45152
rect 9998 45065 10058 45152
rect 10550 45065 10610 45152
rect 11102 45065 11162 45152
rect 11654 45065 11714 45152
rect 12206 45065 12266 45152
rect 12758 45065 12818 45152
rect 13310 45065 13370 45152
rect 13862 45065 13922 45152
rect 14414 45065 14474 45152
rect 14966 45065 15026 45152
rect 15518 45065 15578 45152
rect 16070 45065 16130 45152
rect 16622 45065 16682 45152
rect 17174 45065 17234 45152
rect 17726 45065 17786 45152
rect 18278 45065 18338 45152
rect 18830 45065 18890 45152
rect 6130 44505 6200 45065
rect 6680 44505 6750 45065
rect 7230 44505 7305 45065
rect 7780 44505 7855 45065
rect 8335 44505 8410 45065
rect 8885 44505 8960 45065
rect 9440 44505 9515 45065
rect 9990 44505 10065 45065
rect 10540 44505 10615 45065
rect 11095 44505 11170 45065
rect 11645 44505 11720 45065
rect 12200 44505 12275 45065
rect 12750 44505 12825 45065
rect 13300 44505 13375 45065
rect 13855 44505 13930 45065
rect 14405 44505 14480 45065
rect 14960 44505 15030 45065
rect 15510 44505 15585 45065
rect 16060 44505 16135 45065
rect 16615 44505 16690 45065
rect 17165 44505 17240 45065
rect 17720 44505 17790 45065
rect 18270 44505 18345 45065
rect 18825 44505 18895 45065
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 45060 25514 45152
rect 26006 45060 26066 45152
rect 26558 45060 26618 45152
rect 27110 45060 27170 45152
rect 27662 45060 27722 45152
rect 6130 44280 18895 44505
rect 200 29970 600 44152
rect 200 29645 210 29970
rect 590 29645 600 29970
rect 200 25865 600 29645
rect 200 24700 210 25865
rect 590 24700 600 25865
rect 200 19270 600 24700
rect 200 18945 210 19270
rect 590 18945 600 19270
rect 200 1000 600 18945
rect 800 43645 1200 44152
rect 6130 43645 6355 44280
rect 800 43420 6355 43645
rect 25450 43430 25520 45060
rect 25290 43420 25520 43430
rect 800 40720 1200 43420
rect 25290 43030 25300 43420
rect 25510 43030 25520 43420
rect 25290 43020 25520 43030
rect 26000 40930 26070 45060
rect 26555 41580 26625 45060
rect 27105 42235 27175 45060
rect 27655 42890 27725 45060
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 27655 42880 27820 42890
rect 27655 42780 27665 42880
rect 27810 42780 27820 42880
rect 27655 42770 27820 42780
rect 27105 42225 27270 42235
rect 27105 42125 27115 42225
rect 27260 42125 27270 42225
rect 27105 42115 27270 42125
rect 26555 41570 26720 41580
rect 26555 41470 26565 41570
rect 26710 41470 26720 41570
rect 26555 41460 26720 41470
rect 26000 40920 26165 40930
rect 26000 40820 26010 40920
rect 26155 40820 26165 40920
rect 26000 40810 26165 40820
rect 800 39980 840 40720
rect 1160 39980 1200 40720
rect 800 35580 1200 39980
rect 50135 36630 53280 37250
rect 800 34840 840 35580
rect 1160 34840 1200 35580
rect 800 31635 1200 34840
rect 46965 33335 47585 33885
rect 46965 32715 52290 33335
rect 800 31320 810 31635
rect 1190 31320 1200 31635
rect 800 28800 1200 31320
rect 800 28060 840 28800
rect 1160 28060 1200 28800
rect 51670 28315 52290 32715
rect 52660 31955 53280 36630
rect 52660 31715 52675 31955
rect 53265 31715 53280 31955
rect 52660 31700 53280 31715
rect 51670 28075 51685 28315
rect 52275 28075 52290 28315
rect 51670 28060 52290 28075
rect 800 23215 1200 28060
rect 800 20865 810 23215
rect 1190 20865 1200 23215
rect 800 13860 1200 20865
rect 800 13545 810 13860
rect 1190 13545 1200 13860
rect 800 9320 1200 13545
rect 51670 17615 52290 17630
rect 51670 17375 51685 17615
rect 52275 17375 52290 17615
rect 51670 12565 52290 17375
rect 46735 11945 52290 12565
rect 52660 17085 53280 17100
rect 52660 16845 52675 17085
rect 53265 16845 53280 17085
rect 46735 11395 47355 11945
rect 800 8580 840 9320
rect 1160 8580 1200 9320
rect 52660 8700 53280 16845
rect 800 4120 1200 8580
rect 50140 8080 53280 8700
rect 800 3380 840 4120
rect 1160 3380 1200 4120
rect 26275 4670 26680 4680
rect 26275 4285 26285 4670
rect 26670 4285 26680 4670
rect 800 1000 1200 3380
rect 22410 3615 22815 3625
rect 22410 3230 22420 3615
rect 22805 3230 22815 3615
rect 18545 2545 18950 2555
rect 18545 2160 18555 2545
rect 18940 2160 18950 2545
rect 14680 1505 15085 1515
rect 14680 1140 14690 1505
rect 15075 1140 15085 1505
rect 14680 1130 15085 1140
rect 18545 1130 18950 2160
rect 22410 1130 22815 3230
rect 26275 1130 26680 4285
rect 14905 200 15085 1130
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 1130
rect 22630 200 22815 1130
rect 26495 200 26680 1130
rect 30360 1730 30955 1740
rect 30360 1140 30370 1730
rect 30945 1140 30955 1730
rect 30360 1130 30955 1140
rect 30360 200 30545 1130
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30362 0 30542 200
<< comment >>
rect 63600 44600 66800 45000
rect 66400 400 66800 44600
rect 63600 0 66800 400
use iq_modulator  iq_modulator_0
timestamp 1762794087
transform 1 0 18600 0 1 20200
box -5600 -15200 36430 20020
use sky130_fd_pr__cap_mim_m3_1_DZLWMC  sky130_fd_pr__cap_mim_m3_1_DZLWMC_1
timestamp 1762790939
transform 1 0 47016 0 1 36840
box -3216 -3040 3216 3040
use sky130_fd_pr__cap_mim_m3_1_PP9XRG  sky130_fd_pr__cap_mim_m3_1_PP9XRG_0
timestamp 1762790939
transform 1 0 47016 0 1 8440
box -3216 -3040 3216 3040
use sky130_fd_pr__nfet_01v8_M3JGWT  sky130_fd_pr__nfet_01v8_M3JGWT_0
timestamp 1762799305
transform 1 0 4996 0 1 21973
box -2196 -20973 2196 20973
<< labels >>
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 66976 45152
<< end >>
