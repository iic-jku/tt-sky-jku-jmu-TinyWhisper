magic
tech sky130A
magscale 1 2
timestamp 1762702453
<< metal4 >>
rect -21785 945 395 1050
rect -21785 840 -21680 945
rect -20085 840 -19980 945
rect -18390 840 -18285 945
rect -16690 840 -16585 945
rect -14995 840 -14890 945
rect -13295 840 -13190 945
rect -11600 840 -11495 945
rect -9900 840 -9795 945
rect -8205 840 -8100 945
rect -6505 840 -6400 945
rect -4805 840 -4700 945
rect -3110 840 -3005 945
rect -1410 840 -1305 945
rect 290 840 395 945
rect -21145 -3265 -21040 -3160
rect -19450 -3265 -19345 -3160
rect -17750 -3265 -17645 -3160
rect -16050 -3265 -15945 -3160
rect -14355 -3265 -14250 -3160
rect -12655 -3265 -12550 -3160
rect -10960 -3265 -10855 -3160
rect -9260 -3265 -9155 -3160
rect -7560 -3265 -7455 -3160
rect -5865 -3265 -5760 -3160
rect -4165 -3265 -4060 -3160
rect -2470 -3265 -2365 -3160
rect -770 -3265 -665 -3160
rect 925 -3265 1030 -3160
rect -21145 -3370 1030 -3265
use sky130_fd_pr__cap_mim_m3_1_ZKSXGU  sky130_fd_pr__cap_mim_m3_1_ZKSXGU_0
timestamp 1762702375
transform 1 0 -10521 0 1 -1160
box -11553 -2000 11553 2000
<< labels >>
flabel metal4 -10575 1000 -10575 1000 0 FreeSans 1600 0 0 0 top
port 1 nsew
flabel metal4 -10615 -3320 -10615 -3320 0 FreeSans 1600 0 0 0 bottom
port 3 nsew
<< end >>
