magic
tech sky130A
magscale 1 2
timestamp 1756739912
<< metal3 >>
rect -13251 4312 -12219 4340
rect -13251 3688 -12303 4312
rect -12239 3688 -12219 4312
rect -13251 3660 -12219 3688
rect -11553 4312 -10521 4340
rect -11553 3688 -10605 4312
rect -10541 3688 -10521 4312
rect -11553 3660 -10521 3688
rect -9855 4312 -8823 4340
rect -9855 3688 -8907 4312
rect -8843 3688 -8823 4312
rect -9855 3660 -8823 3688
rect -8157 4312 -7125 4340
rect -8157 3688 -7209 4312
rect -7145 3688 -7125 4312
rect -8157 3660 -7125 3688
rect -6459 4312 -5427 4340
rect -6459 3688 -5511 4312
rect -5447 3688 -5427 4312
rect -6459 3660 -5427 3688
rect -4761 4312 -3729 4340
rect -4761 3688 -3813 4312
rect -3749 3688 -3729 4312
rect -4761 3660 -3729 3688
rect -3063 4312 -2031 4340
rect -3063 3688 -2115 4312
rect -2051 3688 -2031 4312
rect -3063 3660 -2031 3688
rect -1365 4312 -333 4340
rect -1365 3688 -417 4312
rect -353 3688 -333 4312
rect -1365 3660 -333 3688
rect 333 4312 1365 4340
rect 333 3688 1281 4312
rect 1345 3688 1365 4312
rect 333 3660 1365 3688
rect 2031 4312 3063 4340
rect 2031 3688 2979 4312
rect 3043 3688 3063 4312
rect 2031 3660 3063 3688
rect 3729 4312 4761 4340
rect 3729 3688 4677 4312
rect 4741 3688 4761 4312
rect 3729 3660 4761 3688
rect 5427 4312 6459 4340
rect 5427 3688 6375 4312
rect 6439 3688 6459 4312
rect 5427 3660 6459 3688
rect 7125 4312 8157 4340
rect 7125 3688 8073 4312
rect 8137 3688 8157 4312
rect 7125 3660 8157 3688
rect 8823 4312 9855 4340
rect 8823 3688 9771 4312
rect 9835 3688 9855 4312
rect 8823 3660 9855 3688
rect 10521 4312 11553 4340
rect 10521 3688 11469 4312
rect 11533 3688 11553 4312
rect 10521 3660 11553 3688
rect 12219 4312 13251 4340
rect 12219 3688 13167 4312
rect 13231 3688 13251 4312
rect 12219 3660 13251 3688
rect -13251 3312 -12219 3340
rect -13251 2688 -12303 3312
rect -12239 2688 -12219 3312
rect -13251 2660 -12219 2688
rect -11553 3312 -10521 3340
rect -11553 2688 -10605 3312
rect -10541 2688 -10521 3312
rect -11553 2660 -10521 2688
rect -9855 3312 -8823 3340
rect -9855 2688 -8907 3312
rect -8843 2688 -8823 3312
rect -9855 2660 -8823 2688
rect -8157 3312 -7125 3340
rect -8157 2688 -7209 3312
rect -7145 2688 -7125 3312
rect -8157 2660 -7125 2688
rect -6459 3312 -5427 3340
rect -6459 2688 -5511 3312
rect -5447 2688 -5427 3312
rect -6459 2660 -5427 2688
rect -4761 3312 -3729 3340
rect -4761 2688 -3813 3312
rect -3749 2688 -3729 3312
rect -4761 2660 -3729 2688
rect -3063 3312 -2031 3340
rect -3063 2688 -2115 3312
rect -2051 2688 -2031 3312
rect -3063 2660 -2031 2688
rect -1365 3312 -333 3340
rect -1365 2688 -417 3312
rect -353 2688 -333 3312
rect -1365 2660 -333 2688
rect 333 3312 1365 3340
rect 333 2688 1281 3312
rect 1345 2688 1365 3312
rect 333 2660 1365 2688
rect 2031 3312 3063 3340
rect 2031 2688 2979 3312
rect 3043 2688 3063 3312
rect 2031 2660 3063 2688
rect 3729 3312 4761 3340
rect 3729 2688 4677 3312
rect 4741 2688 4761 3312
rect 3729 2660 4761 2688
rect 5427 3312 6459 3340
rect 5427 2688 6375 3312
rect 6439 2688 6459 3312
rect 5427 2660 6459 2688
rect 7125 3312 8157 3340
rect 7125 2688 8073 3312
rect 8137 2688 8157 3312
rect 7125 2660 8157 2688
rect 8823 3312 9855 3340
rect 8823 2688 9771 3312
rect 9835 2688 9855 3312
rect 8823 2660 9855 2688
rect 10521 3312 11553 3340
rect 10521 2688 11469 3312
rect 11533 2688 11553 3312
rect 10521 2660 11553 2688
rect 12219 3312 13251 3340
rect 12219 2688 13167 3312
rect 13231 2688 13251 3312
rect 12219 2660 13251 2688
rect -13251 2312 -12219 2340
rect -13251 1688 -12303 2312
rect -12239 1688 -12219 2312
rect -13251 1660 -12219 1688
rect -11553 2312 -10521 2340
rect -11553 1688 -10605 2312
rect -10541 1688 -10521 2312
rect -11553 1660 -10521 1688
rect -9855 2312 -8823 2340
rect -9855 1688 -8907 2312
rect -8843 1688 -8823 2312
rect -9855 1660 -8823 1688
rect -8157 2312 -7125 2340
rect -8157 1688 -7209 2312
rect -7145 1688 -7125 2312
rect -8157 1660 -7125 1688
rect -6459 2312 -5427 2340
rect -6459 1688 -5511 2312
rect -5447 1688 -5427 2312
rect -6459 1660 -5427 1688
rect -4761 2312 -3729 2340
rect -4761 1688 -3813 2312
rect -3749 1688 -3729 2312
rect -4761 1660 -3729 1688
rect -3063 2312 -2031 2340
rect -3063 1688 -2115 2312
rect -2051 1688 -2031 2312
rect -3063 1660 -2031 1688
rect -1365 2312 -333 2340
rect -1365 1688 -417 2312
rect -353 1688 -333 2312
rect -1365 1660 -333 1688
rect 333 2312 1365 2340
rect 333 1688 1281 2312
rect 1345 1688 1365 2312
rect 333 1660 1365 1688
rect 2031 2312 3063 2340
rect 2031 1688 2979 2312
rect 3043 1688 3063 2312
rect 2031 1660 3063 1688
rect 3729 2312 4761 2340
rect 3729 1688 4677 2312
rect 4741 1688 4761 2312
rect 3729 1660 4761 1688
rect 5427 2312 6459 2340
rect 5427 1688 6375 2312
rect 6439 1688 6459 2312
rect 5427 1660 6459 1688
rect 7125 2312 8157 2340
rect 7125 1688 8073 2312
rect 8137 1688 8157 2312
rect 7125 1660 8157 1688
rect 8823 2312 9855 2340
rect 8823 1688 9771 2312
rect 9835 1688 9855 2312
rect 8823 1660 9855 1688
rect 10521 2312 11553 2340
rect 10521 1688 11469 2312
rect 11533 1688 11553 2312
rect 10521 1660 11553 1688
rect 12219 2312 13251 2340
rect 12219 1688 13167 2312
rect 13231 1688 13251 2312
rect 12219 1660 13251 1688
rect -13251 1312 -12219 1340
rect -13251 688 -12303 1312
rect -12239 688 -12219 1312
rect -13251 660 -12219 688
rect -11553 1312 -10521 1340
rect -11553 688 -10605 1312
rect -10541 688 -10521 1312
rect -11553 660 -10521 688
rect -9855 1312 -8823 1340
rect -9855 688 -8907 1312
rect -8843 688 -8823 1312
rect -9855 660 -8823 688
rect -8157 1312 -7125 1340
rect -8157 688 -7209 1312
rect -7145 688 -7125 1312
rect -8157 660 -7125 688
rect -6459 1312 -5427 1340
rect -6459 688 -5511 1312
rect -5447 688 -5427 1312
rect -6459 660 -5427 688
rect -4761 1312 -3729 1340
rect -4761 688 -3813 1312
rect -3749 688 -3729 1312
rect -4761 660 -3729 688
rect -3063 1312 -2031 1340
rect -3063 688 -2115 1312
rect -2051 688 -2031 1312
rect -3063 660 -2031 688
rect -1365 1312 -333 1340
rect -1365 688 -417 1312
rect -353 688 -333 1312
rect -1365 660 -333 688
rect 333 1312 1365 1340
rect 333 688 1281 1312
rect 1345 688 1365 1312
rect 333 660 1365 688
rect 2031 1312 3063 1340
rect 2031 688 2979 1312
rect 3043 688 3063 1312
rect 2031 660 3063 688
rect 3729 1312 4761 1340
rect 3729 688 4677 1312
rect 4741 688 4761 1312
rect 3729 660 4761 688
rect 5427 1312 6459 1340
rect 5427 688 6375 1312
rect 6439 688 6459 1312
rect 5427 660 6459 688
rect 7125 1312 8157 1340
rect 7125 688 8073 1312
rect 8137 688 8157 1312
rect 7125 660 8157 688
rect 8823 1312 9855 1340
rect 8823 688 9771 1312
rect 9835 688 9855 1312
rect 8823 660 9855 688
rect 10521 1312 11553 1340
rect 10521 688 11469 1312
rect 11533 688 11553 1312
rect 10521 660 11553 688
rect 12219 1312 13251 1340
rect 12219 688 13167 1312
rect 13231 688 13251 1312
rect 12219 660 13251 688
rect -13251 312 -12219 340
rect -13251 -312 -12303 312
rect -12239 -312 -12219 312
rect -13251 -340 -12219 -312
rect -11553 312 -10521 340
rect -11553 -312 -10605 312
rect -10541 -312 -10521 312
rect -11553 -340 -10521 -312
rect -9855 312 -8823 340
rect -9855 -312 -8907 312
rect -8843 -312 -8823 312
rect -9855 -340 -8823 -312
rect -8157 312 -7125 340
rect -8157 -312 -7209 312
rect -7145 -312 -7125 312
rect -8157 -340 -7125 -312
rect -6459 312 -5427 340
rect -6459 -312 -5511 312
rect -5447 -312 -5427 312
rect -6459 -340 -5427 -312
rect -4761 312 -3729 340
rect -4761 -312 -3813 312
rect -3749 -312 -3729 312
rect -4761 -340 -3729 -312
rect -3063 312 -2031 340
rect -3063 -312 -2115 312
rect -2051 -312 -2031 312
rect -3063 -340 -2031 -312
rect -1365 312 -333 340
rect -1365 -312 -417 312
rect -353 -312 -333 312
rect -1365 -340 -333 -312
rect 333 312 1365 340
rect 333 -312 1281 312
rect 1345 -312 1365 312
rect 333 -340 1365 -312
rect 2031 312 3063 340
rect 2031 -312 2979 312
rect 3043 -312 3063 312
rect 2031 -340 3063 -312
rect 3729 312 4761 340
rect 3729 -312 4677 312
rect 4741 -312 4761 312
rect 3729 -340 4761 -312
rect 5427 312 6459 340
rect 5427 -312 6375 312
rect 6439 -312 6459 312
rect 5427 -340 6459 -312
rect 7125 312 8157 340
rect 7125 -312 8073 312
rect 8137 -312 8157 312
rect 7125 -340 8157 -312
rect 8823 312 9855 340
rect 8823 -312 9771 312
rect 9835 -312 9855 312
rect 8823 -340 9855 -312
rect 10521 312 11553 340
rect 10521 -312 11469 312
rect 11533 -312 11553 312
rect 10521 -340 11553 -312
rect 12219 312 13251 340
rect 12219 -312 13167 312
rect 13231 -312 13251 312
rect 12219 -340 13251 -312
rect -13251 -688 -12219 -660
rect -13251 -1312 -12303 -688
rect -12239 -1312 -12219 -688
rect -13251 -1340 -12219 -1312
rect -11553 -688 -10521 -660
rect -11553 -1312 -10605 -688
rect -10541 -1312 -10521 -688
rect -11553 -1340 -10521 -1312
rect -9855 -688 -8823 -660
rect -9855 -1312 -8907 -688
rect -8843 -1312 -8823 -688
rect -9855 -1340 -8823 -1312
rect -8157 -688 -7125 -660
rect -8157 -1312 -7209 -688
rect -7145 -1312 -7125 -688
rect -8157 -1340 -7125 -1312
rect -6459 -688 -5427 -660
rect -6459 -1312 -5511 -688
rect -5447 -1312 -5427 -688
rect -6459 -1340 -5427 -1312
rect -4761 -688 -3729 -660
rect -4761 -1312 -3813 -688
rect -3749 -1312 -3729 -688
rect -4761 -1340 -3729 -1312
rect -3063 -688 -2031 -660
rect -3063 -1312 -2115 -688
rect -2051 -1312 -2031 -688
rect -3063 -1340 -2031 -1312
rect -1365 -688 -333 -660
rect -1365 -1312 -417 -688
rect -353 -1312 -333 -688
rect -1365 -1340 -333 -1312
rect 333 -688 1365 -660
rect 333 -1312 1281 -688
rect 1345 -1312 1365 -688
rect 333 -1340 1365 -1312
rect 2031 -688 3063 -660
rect 2031 -1312 2979 -688
rect 3043 -1312 3063 -688
rect 2031 -1340 3063 -1312
rect 3729 -688 4761 -660
rect 3729 -1312 4677 -688
rect 4741 -1312 4761 -688
rect 3729 -1340 4761 -1312
rect 5427 -688 6459 -660
rect 5427 -1312 6375 -688
rect 6439 -1312 6459 -688
rect 5427 -1340 6459 -1312
rect 7125 -688 8157 -660
rect 7125 -1312 8073 -688
rect 8137 -1312 8157 -688
rect 7125 -1340 8157 -1312
rect 8823 -688 9855 -660
rect 8823 -1312 9771 -688
rect 9835 -1312 9855 -688
rect 8823 -1340 9855 -1312
rect 10521 -688 11553 -660
rect 10521 -1312 11469 -688
rect 11533 -1312 11553 -688
rect 10521 -1340 11553 -1312
rect 12219 -688 13251 -660
rect 12219 -1312 13167 -688
rect 13231 -1312 13251 -688
rect 12219 -1340 13251 -1312
rect -13251 -1688 -12219 -1660
rect -13251 -2312 -12303 -1688
rect -12239 -2312 -12219 -1688
rect -13251 -2340 -12219 -2312
rect -11553 -1688 -10521 -1660
rect -11553 -2312 -10605 -1688
rect -10541 -2312 -10521 -1688
rect -11553 -2340 -10521 -2312
rect -9855 -1688 -8823 -1660
rect -9855 -2312 -8907 -1688
rect -8843 -2312 -8823 -1688
rect -9855 -2340 -8823 -2312
rect -8157 -1688 -7125 -1660
rect -8157 -2312 -7209 -1688
rect -7145 -2312 -7125 -1688
rect -8157 -2340 -7125 -2312
rect -6459 -1688 -5427 -1660
rect -6459 -2312 -5511 -1688
rect -5447 -2312 -5427 -1688
rect -6459 -2340 -5427 -2312
rect -4761 -1688 -3729 -1660
rect -4761 -2312 -3813 -1688
rect -3749 -2312 -3729 -1688
rect -4761 -2340 -3729 -2312
rect -3063 -1688 -2031 -1660
rect -3063 -2312 -2115 -1688
rect -2051 -2312 -2031 -1688
rect -3063 -2340 -2031 -2312
rect -1365 -1688 -333 -1660
rect -1365 -2312 -417 -1688
rect -353 -2312 -333 -1688
rect -1365 -2340 -333 -2312
rect 333 -1688 1365 -1660
rect 333 -2312 1281 -1688
rect 1345 -2312 1365 -1688
rect 333 -2340 1365 -2312
rect 2031 -1688 3063 -1660
rect 2031 -2312 2979 -1688
rect 3043 -2312 3063 -1688
rect 2031 -2340 3063 -2312
rect 3729 -1688 4761 -1660
rect 3729 -2312 4677 -1688
rect 4741 -2312 4761 -1688
rect 3729 -2340 4761 -2312
rect 5427 -1688 6459 -1660
rect 5427 -2312 6375 -1688
rect 6439 -2312 6459 -1688
rect 5427 -2340 6459 -2312
rect 7125 -1688 8157 -1660
rect 7125 -2312 8073 -1688
rect 8137 -2312 8157 -1688
rect 7125 -2340 8157 -2312
rect 8823 -1688 9855 -1660
rect 8823 -2312 9771 -1688
rect 9835 -2312 9855 -1688
rect 8823 -2340 9855 -2312
rect 10521 -1688 11553 -1660
rect 10521 -2312 11469 -1688
rect 11533 -2312 11553 -1688
rect 10521 -2340 11553 -2312
rect 12219 -1688 13251 -1660
rect 12219 -2312 13167 -1688
rect 13231 -2312 13251 -1688
rect 12219 -2340 13251 -2312
rect -13251 -2688 -12219 -2660
rect -13251 -3312 -12303 -2688
rect -12239 -3312 -12219 -2688
rect -13251 -3340 -12219 -3312
rect -11553 -2688 -10521 -2660
rect -11553 -3312 -10605 -2688
rect -10541 -3312 -10521 -2688
rect -11553 -3340 -10521 -3312
rect -9855 -2688 -8823 -2660
rect -9855 -3312 -8907 -2688
rect -8843 -3312 -8823 -2688
rect -9855 -3340 -8823 -3312
rect -8157 -2688 -7125 -2660
rect -8157 -3312 -7209 -2688
rect -7145 -3312 -7125 -2688
rect -8157 -3340 -7125 -3312
rect -6459 -2688 -5427 -2660
rect -6459 -3312 -5511 -2688
rect -5447 -3312 -5427 -2688
rect -6459 -3340 -5427 -3312
rect -4761 -2688 -3729 -2660
rect -4761 -3312 -3813 -2688
rect -3749 -3312 -3729 -2688
rect -4761 -3340 -3729 -3312
rect -3063 -2688 -2031 -2660
rect -3063 -3312 -2115 -2688
rect -2051 -3312 -2031 -2688
rect -3063 -3340 -2031 -3312
rect -1365 -2688 -333 -2660
rect -1365 -3312 -417 -2688
rect -353 -3312 -333 -2688
rect -1365 -3340 -333 -3312
rect 333 -2688 1365 -2660
rect 333 -3312 1281 -2688
rect 1345 -3312 1365 -2688
rect 333 -3340 1365 -3312
rect 2031 -2688 3063 -2660
rect 2031 -3312 2979 -2688
rect 3043 -3312 3063 -2688
rect 2031 -3340 3063 -3312
rect 3729 -2688 4761 -2660
rect 3729 -3312 4677 -2688
rect 4741 -3312 4761 -2688
rect 3729 -3340 4761 -3312
rect 5427 -2688 6459 -2660
rect 5427 -3312 6375 -2688
rect 6439 -3312 6459 -2688
rect 5427 -3340 6459 -3312
rect 7125 -2688 8157 -2660
rect 7125 -3312 8073 -2688
rect 8137 -3312 8157 -2688
rect 7125 -3340 8157 -3312
rect 8823 -2688 9855 -2660
rect 8823 -3312 9771 -2688
rect 9835 -3312 9855 -2688
rect 8823 -3340 9855 -3312
rect 10521 -2688 11553 -2660
rect 10521 -3312 11469 -2688
rect 11533 -3312 11553 -2688
rect 10521 -3340 11553 -3312
rect 12219 -2688 13251 -2660
rect 12219 -3312 13167 -2688
rect 13231 -3312 13251 -2688
rect 12219 -3340 13251 -3312
rect -13251 -3688 -12219 -3660
rect -13251 -4312 -12303 -3688
rect -12239 -4312 -12219 -3688
rect -13251 -4340 -12219 -4312
rect -11553 -3688 -10521 -3660
rect -11553 -4312 -10605 -3688
rect -10541 -4312 -10521 -3688
rect -11553 -4340 -10521 -4312
rect -9855 -3688 -8823 -3660
rect -9855 -4312 -8907 -3688
rect -8843 -4312 -8823 -3688
rect -9855 -4340 -8823 -4312
rect -8157 -3688 -7125 -3660
rect -8157 -4312 -7209 -3688
rect -7145 -4312 -7125 -3688
rect -8157 -4340 -7125 -4312
rect -6459 -3688 -5427 -3660
rect -6459 -4312 -5511 -3688
rect -5447 -4312 -5427 -3688
rect -6459 -4340 -5427 -4312
rect -4761 -3688 -3729 -3660
rect -4761 -4312 -3813 -3688
rect -3749 -4312 -3729 -3688
rect -4761 -4340 -3729 -4312
rect -3063 -3688 -2031 -3660
rect -3063 -4312 -2115 -3688
rect -2051 -4312 -2031 -3688
rect -3063 -4340 -2031 -4312
rect -1365 -3688 -333 -3660
rect -1365 -4312 -417 -3688
rect -353 -4312 -333 -3688
rect -1365 -4340 -333 -4312
rect 333 -3688 1365 -3660
rect 333 -4312 1281 -3688
rect 1345 -4312 1365 -3688
rect 333 -4340 1365 -4312
rect 2031 -3688 3063 -3660
rect 2031 -4312 2979 -3688
rect 3043 -4312 3063 -3688
rect 2031 -4340 3063 -4312
rect 3729 -3688 4761 -3660
rect 3729 -4312 4677 -3688
rect 4741 -4312 4761 -3688
rect 3729 -4340 4761 -4312
rect 5427 -3688 6459 -3660
rect 5427 -4312 6375 -3688
rect 6439 -4312 6459 -3688
rect 5427 -4340 6459 -4312
rect 7125 -3688 8157 -3660
rect 7125 -4312 8073 -3688
rect 8137 -4312 8157 -3688
rect 7125 -4340 8157 -4312
rect 8823 -3688 9855 -3660
rect 8823 -4312 9771 -3688
rect 9835 -4312 9855 -3688
rect 8823 -4340 9855 -4312
rect 10521 -3688 11553 -3660
rect 10521 -4312 11469 -3688
rect 11533 -4312 11553 -3688
rect 10521 -4340 11553 -4312
rect 12219 -3688 13251 -3660
rect 12219 -4312 13167 -3688
rect 13231 -4312 13251 -3688
rect 12219 -4340 13251 -4312
<< via3 >>
rect -12303 3688 -12239 4312
rect -10605 3688 -10541 4312
rect -8907 3688 -8843 4312
rect -7209 3688 -7145 4312
rect -5511 3688 -5447 4312
rect -3813 3688 -3749 4312
rect -2115 3688 -2051 4312
rect -417 3688 -353 4312
rect 1281 3688 1345 4312
rect 2979 3688 3043 4312
rect 4677 3688 4741 4312
rect 6375 3688 6439 4312
rect 8073 3688 8137 4312
rect 9771 3688 9835 4312
rect 11469 3688 11533 4312
rect 13167 3688 13231 4312
rect -12303 2688 -12239 3312
rect -10605 2688 -10541 3312
rect -8907 2688 -8843 3312
rect -7209 2688 -7145 3312
rect -5511 2688 -5447 3312
rect -3813 2688 -3749 3312
rect -2115 2688 -2051 3312
rect -417 2688 -353 3312
rect 1281 2688 1345 3312
rect 2979 2688 3043 3312
rect 4677 2688 4741 3312
rect 6375 2688 6439 3312
rect 8073 2688 8137 3312
rect 9771 2688 9835 3312
rect 11469 2688 11533 3312
rect 13167 2688 13231 3312
rect -12303 1688 -12239 2312
rect -10605 1688 -10541 2312
rect -8907 1688 -8843 2312
rect -7209 1688 -7145 2312
rect -5511 1688 -5447 2312
rect -3813 1688 -3749 2312
rect -2115 1688 -2051 2312
rect -417 1688 -353 2312
rect 1281 1688 1345 2312
rect 2979 1688 3043 2312
rect 4677 1688 4741 2312
rect 6375 1688 6439 2312
rect 8073 1688 8137 2312
rect 9771 1688 9835 2312
rect 11469 1688 11533 2312
rect 13167 1688 13231 2312
rect -12303 688 -12239 1312
rect -10605 688 -10541 1312
rect -8907 688 -8843 1312
rect -7209 688 -7145 1312
rect -5511 688 -5447 1312
rect -3813 688 -3749 1312
rect -2115 688 -2051 1312
rect -417 688 -353 1312
rect 1281 688 1345 1312
rect 2979 688 3043 1312
rect 4677 688 4741 1312
rect 6375 688 6439 1312
rect 8073 688 8137 1312
rect 9771 688 9835 1312
rect 11469 688 11533 1312
rect 13167 688 13231 1312
rect -12303 -312 -12239 312
rect -10605 -312 -10541 312
rect -8907 -312 -8843 312
rect -7209 -312 -7145 312
rect -5511 -312 -5447 312
rect -3813 -312 -3749 312
rect -2115 -312 -2051 312
rect -417 -312 -353 312
rect 1281 -312 1345 312
rect 2979 -312 3043 312
rect 4677 -312 4741 312
rect 6375 -312 6439 312
rect 8073 -312 8137 312
rect 9771 -312 9835 312
rect 11469 -312 11533 312
rect 13167 -312 13231 312
rect -12303 -1312 -12239 -688
rect -10605 -1312 -10541 -688
rect -8907 -1312 -8843 -688
rect -7209 -1312 -7145 -688
rect -5511 -1312 -5447 -688
rect -3813 -1312 -3749 -688
rect -2115 -1312 -2051 -688
rect -417 -1312 -353 -688
rect 1281 -1312 1345 -688
rect 2979 -1312 3043 -688
rect 4677 -1312 4741 -688
rect 6375 -1312 6439 -688
rect 8073 -1312 8137 -688
rect 9771 -1312 9835 -688
rect 11469 -1312 11533 -688
rect 13167 -1312 13231 -688
rect -12303 -2312 -12239 -1688
rect -10605 -2312 -10541 -1688
rect -8907 -2312 -8843 -1688
rect -7209 -2312 -7145 -1688
rect -5511 -2312 -5447 -1688
rect -3813 -2312 -3749 -1688
rect -2115 -2312 -2051 -1688
rect -417 -2312 -353 -1688
rect 1281 -2312 1345 -1688
rect 2979 -2312 3043 -1688
rect 4677 -2312 4741 -1688
rect 6375 -2312 6439 -1688
rect 8073 -2312 8137 -1688
rect 9771 -2312 9835 -1688
rect 11469 -2312 11533 -1688
rect 13167 -2312 13231 -1688
rect -12303 -3312 -12239 -2688
rect -10605 -3312 -10541 -2688
rect -8907 -3312 -8843 -2688
rect -7209 -3312 -7145 -2688
rect -5511 -3312 -5447 -2688
rect -3813 -3312 -3749 -2688
rect -2115 -3312 -2051 -2688
rect -417 -3312 -353 -2688
rect 1281 -3312 1345 -2688
rect 2979 -3312 3043 -2688
rect 4677 -3312 4741 -2688
rect 6375 -3312 6439 -2688
rect 8073 -3312 8137 -2688
rect 9771 -3312 9835 -2688
rect 11469 -3312 11533 -2688
rect 13167 -3312 13231 -2688
rect -12303 -4312 -12239 -3688
rect -10605 -4312 -10541 -3688
rect -8907 -4312 -8843 -3688
rect -7209 -4312 -7145 -3688
rect -5511 -4312 -5447 -3688
rect -3813 -4312 -3749 -3688
rect -2115 -4312 -2051 -3688
rect -417 -4312 -353 -3688
rect 1281 -4312 1345 -3688
rect 2979 -4312 3043 -3688
rect 4677 -4312 4741 -3688
rect 6375 -4312 6439 -3688
rect 8073 -4312 8137 -3688
rect 9771 -4312 9835 -3688
rect 11469 -4312 11533 -3688
rect 13167 -4312 13231 -3688
<< mimcap >>
rect -13211 4260 -12611 4300
rect -13211 3740 -13171 4260
rect -12651 3740 -12611 4260
rect -13211 3700 -12611 3740
rect -11513 4260 -10913 4300
rect -11513 3740 -11473 4260
rect -10953 3740 -10913 4260
rect -11513 3700 -10913 3740
rect -9815 4260 -9215 4300
rect -9815 3740 -9775 4260
rect -9255 3740 -9215 4260
rect -9815 3700 -9215 3740
rect -8117 4260 -7517 4300
rect -8117 3740 -8077 4260
rect -7557 3740 -7517 4260
rect -8117 3700 -7517 3740
rect -6419 4260 -5819 4300
rect -6419 3740 -6379 4260
rect -5859 3740 -5819 4260
rect -6419 3700 -5819 3740
rect -4721 4260 -4121 4300
rect -4721 3740 -4681 4260
rect -4161 3740 -4121 4260
rect -4721 3700 -4121 3740
rect -3023 4260 -2423 4300
rect -3023 3740 -2983 4260
rect -2463 3740 -2423 4260
rect -3023 3700 -2423 3740
rect -1325 4260 -725 4300
rect -1325 3740 -1285 4260
rect -765 3740 -725 4260
rect -1325 3700 -725 3740
rect 373 4260 973 4300
rect 373 3740 413 4260
rect 933 3740 973 4260
rect 373 3700 973 3740
rect 2071 4260 2671 4300
rect 2071 3740 2111 4260
rect 2631 3740 2671 4260
rect 2071 3700 2671 3740
rect 3769 4260 4369 4300
rect 3769 3740 3809 4260
rect 4329 3740 4369 4260
rect 3769 3700 4369 3740
rect 5467 4260 6067 4300
rect 5467 3740 5507 4260
rect 6027 3740 6067 4260
rect 5467 3700 6067 3740
rect 7165 4260 7765 4300
rect 7165 3740 7205 4260
rect 7725 3740 7765 4260
rect 7165 3700 7765 3740
rect 8863 4260 9463 4300
rect 8863 3740 8903 4260
rect 9423 3740 9463 4260
rect 8863 3700 9463 3740
rect 10561 4260 11161 4300
rect 10561 3740 10601 4260
rect 11121 3740 11161 4260
rect 10561 3700 11161 3740
rect 12259 4260 12859 4300
rect 12259 3740 12299 4260
rect 12819 3740 12859 4260
rect 12259 3700 12859 3740
rect -13211 3260 -12611 3300
rect -13211 2740 -13171 3260
rect -12651 2740 -12611 3260
rect -13211 2700 -12611 2740
rect -11513 3260 -10913 3300
rect -11513 2740 -11473 3260
rect -10953 2740 -10913 3260
rect -11513 2700 -10913 2740
rect -9815 3260 -9215 3300
rect -9815 2740 -9775 3260
rect -9255 2740 -9215 3260
rect -9815 2700 -9215 2740
rect -8117 3260 -7517 3300
rect -8117 2740 -8077 3260
rect -7557 2740 -7517 3260
rect -8117 2700 -7517 2740
rect -6419 3260 -5819 3300
rect -6419 2740 -6379 3260
rect -5859 2740 -5819 3260
rect -6419 2700 -5819 2740
rect -4721 3260 -4121 3300
rect -4721 2740 -4681 3260
rect -4161 2740 -4121 3260
rect -4721 2700 -4121 2740
rect -3023 3260 -2423 3300
rect -3023 2740 -2983 3260
rect -2463 2740 -2423 3260
rect -3023 2700 -2423 2740
rect -1325 3260 -725 3300
rect -1325 2740 -1285 3260
rect -765 2740 -725 3260
rect -1325 2700 -725 2740
rect 373 3260 973 3300
rect 373 2740 413 3260
rect 933 2740 973 3260
rect 373 2700 973 2740
rect 2071 3260 2671 3300
rect 2071 2740 2111 3260
rect 2631 2740 2671 3260
rect 2071 2700 2671 2740
rect 3769 3260 4369 3300
rect 3769 2740 3809 3260
rect 4329 2740 4369 3260
rect 3769 2700 4369 2740
rect 5467 3260 6067 3300
rect 5467 2740 5507 3260
rect 6027 2740 6067 3260
rect 5467 2700 6067 2740
rect 7165 3260 7765 3300
rect 7165 2740 7205 3260
rect 7725 2740 7765 3260
rect 7165 2700 7765 2740
rect 8863 3260 9463 3300
rect 8863 2740 8903 3260
rect 9423 2740 9463 3260
rect 8863 2700 9463 2740
rect 10561 3260 11161 3300
rect 10561 2740 10601 3260
rect 11121 2740 11161 3260
rect 10561 2700 11161 2740
rect 12259 3260 12859 3300
rect 12259 2740 12299 3260
rect 12819 2740 12859 3260
rect 12259 2700 12859 2740
rect -13211 2260 -12611 2300
rect -13211 1740 -13171 2260
rect -12651 1740 -12611 2260
rect -13211 1700 -12611 1740
rect -11513 2260 -10913 2300
rect -11513 1740 -11473 2260
rect -10953 1740 -10913 2260
rect -11513 1700 -10913 1740
rect -9815 2260 -9215 2300
rect -9815 1740 -9775 2260
rect -9255 1740 -9215 2260
rect -9815 1700 -9215 1740
rect -8117 2260 -7517 2300
rect -8117 1740 -8077 2260
rect -7557 1740 -7517 2260
rect -8117 1700 -7517 1740
rect -6419 2260 -5819 2300
rect -6419 1740 -6379 2260
rect -5859 1740 -5819 2260
rect -6419 1700 -5819 1740
rect -4721 2260 -4121 2300
rect -4721 1740 -4681 2260
rect -4161 1740 -4121 2260
rect -4721 1700 -4121 1740
rect -3023 2260 -2423 2300
rect -3023 1740 -2983 2260
rect -2463 1740 -2423 2260
rect -3023 1700 -2423 1740
rect -1325 2260 -725 2300
rect -1325 1740 -1285 2260
rect -765 1740 -725 2260
rect -1325 1700 -725 1740
rect 373 2260 973 2300
rect 373 1740 413 2260
rect 933 1740 973 2260
rect 373 1700 973 1740
rect 2071 2260 2671 2300
rect 2071 1740 2111 2260
rect 2631 1740 2671 2260
rect 2071 1700 2671 1740
rect 3769 2260 4369 2300
rect 3769 1740 3809 2260
rect 4329 1740 4369 2260
rect 3769 1700 4369 1740
rect 5467 2260 6067 2300
rect 5467 1740 5507 2260
rect 6027 1740 6067 2260
rect 5467 1700 6067 1740
rect 7165 2260 7765 2300
rect 7165 1740 7205 2260
rect 7725 1740 7765 2260
rect 7165 1700 7765 1740
rect 8863 2260 9463 2300
rect 8863 1740 8903 2260
rect 9423 1740 9463 2260
rect 8863 1700 9463 1740
rect 10561 2260 11161 2300
rect 10561 1740 10601 2260
rect 11121 1740 11161 2260
rect 10561 1700 11161 1740
rect 12259 2260 12859 2300
rect 12259 1740 12299 2260
rect 12819 1740 12859 2260
rect 12259 1700 12859 1740
rect -13211 1260 -12611 1300
rect -13211 740 -13171 1260
rect -12651 740 -12611 1260
rect -13211 700 -12611 740
rect -11513 1260 -10913 1300
rect -11513 740 -11473 1260
rect -10953 740 -10913 1260
rect -11513 700 -10913 740
rect -9815 1260 -9215 1300
rect -9815 740 -9775 1260
rect -9255 740 -9215 1260
rect -9815 700 -9215 740
rect -8117 1260 -7517 1300
rect -8117 740 -8077 1260
rect -7557 740 -7517 1260
rect -8117 700 -7517 740
rect -6419 1260 -5819 1300
rect -6419 740 -6379 1260
rect -5859 740 -5819 1260
rect -6419 700 -5819 740
rect -4721 1260 -4121 1300
rect -4721 740 -4681 1260
rect -4161 740 -4121 1260
rect -4721 700 -4121 740
rect -3023 1260 -2423 1300
rect -3023 740 -2983 1260
rect -2463 740 -2423 1260
rect -3023 700 -2423 740
rect -1325 1260 -725 1300
rect -1325 740 -1285 1260
rect -765 740 -725 1260
rect -1325 700 -725 740
rect 373 1260 973 1300
rect 373 740 413 1260
rect 933 740 973 1260
rect 373 700 973 740
rect 2071 1260 2671 1300
rect 2071 740 2111 1260
rect 2631 740 2671 1260
rect 2071 700 2671 740
rect 3769 1260 4369 1300
rect 3769 740 3809 1260
rect 4329 740 4369 1260
rect 3769 700 4369 740
rect 5467 1260 6067 1300
rect 5467 740 5507 1260
rect 6027 740 6067 1260
rect 5467 700 6067 740
rect 7165 1260 7765 1300
rect 7165 740 7205 1260
rect 7725 740 7765 1260
rect 7165 700 7765 740
rect 8863 1260 9463 1300
rect 8863 740 8903 1260
rect 9423 740 9463 1260
rect 8863 700 9463 740
rect 10561 1260 11161 1300
rect 10561 740 10601 1260
rect 11121 740 11161 1260
rect 10561 700 11161 740
rect 12259 1260 12859 1300
rect 12259 740 12299 1260
rect 12819 740 12859 1260
rect 12259 700 12859 740
rect -13211 260 -12611 300
rect -13211 -260 -13171 260
rect -12651 -260 -12611 260
rect -13211 -300 -12611 -260
rect -11513 260 -10913 300
rect -11513 -260 -11473 260
rect -10953 -260 -10913 260
rect -11513 -300 -10913 -260
rect -9815 260 -9215 300
rect -9815 -260 -9775 260
rect -9255 -260 -9215 260
rect -9815 -300 -9215 -260
rect -8117 260 -7517 300
rect -8117 -260 -8077 260
rect -7557 -260 -7517 260
rect -8117 -300 -7517 -260
rect -6419 260 -5819 300
rect -6419 -260 -6379 260
rect -5859 -260 -5819 260
rect -6419 -300 -5819 -260
rect -4721 260 -4121 300
rect -4721 -260 -4681 260
rect -4161 -260 -4121 260
rect -4721 -300 -4121 -260
rect -3023 260 -2423 300
rect -3023 -260 -2983 260
rect -2463 -260 -2423 260
rect -3023 -300 -2423 -260
rect -1325 260 -725 300
rect -1325 -260 -1285 260
rect -765 -260 -725 260
rect -1325 -300 -725 -260
rect 373 260 973 300
rect 373 -260 413 260
rect 933 -260 973 260
rect 373 -300 973 -260
rect 2071 260 2671 300
rect 2071 -260 2111 260
rect 2631 -260 2671 260
rect 2071 -300 2671 -260
rect 3769 260 4369 300
rect 3769 -260 3809 260
rect 4329 -260 4369 260
rect 3769 -300 4369 -260
rect 5467 260 6067 300
rect 5467 -260 5507 260
rect 6027 -260 6067 260
rect 5467 -300 6067 -260
rect 7165 260 7765 300
rect 7165 -260 7205 260
rect 7725 -260 7765 260
rect 7165 -300 7765 -260
rect 8863 260 9463 300
rect 8863 -260 8903 260
rect 9423 -260 9463 260
rect 8863 -300 9463 -260
rect 10561 260 11161 300
rect 10561 -260 10601 260
rect 11121 -260 11161 260
rect 10561 -300 11161 -260
rect 12259 260 12859 300
rect 12259 -260 12299 260
rect 12819 -260 12859 260
rect 12259 -300 12859 -260
rect -13211 -740 -12611 -700
rect -13211 -1260 -13171 -740
rect -12651 -1260 -12611 -740
rect -13211 -1300 -12611 -1260
rect -11513 -740 -10913 -700
rect -11513 -1260 -11473 -740
rect -10953 -1260 -10913 -740
rect -11513 -1300 -10913 -1260
rect -9815 -740 -9215 -700
rect -9815 -1260 -9775 -740
rect -9255 -1260 -9215 -740
rect -9815 -1300 -9215 -1260
rect -8117 -740 -7517 -700
rect -8117 -1260 -8077 -740
rect -7557 -1260 -7517 -740
rect -8117 -1300 -7517 -1260
rect -6419 -740 -5819 -700
rect -6419 -1260 -6379 -740
rect -5859 -1260 -5819 -740
rect -6419 -1300 -5819 -1260
rect -4721 -740 -4121 -700
rect -4721 -1260 -4681 -740
rect -4161 -1260 -4121 -740
rect -4721 -1300 -4121 -1260
rect -3023 -740 -2423 -700
rect -3023 -1260 -2983 -740
rect -2463 -1260 -2423 -740
rect -3023 -1300 -2423 -1260
rect -1325 -740 -725 -700
rect -1325 -1260 -1285 -740
rect -765 -1260 -725 -740
rect -1325 -1300 -725 -1260
rect 373 -740 973 -700
rect 373 -1260 413 -740
rect 933 -1260 973 -740
rect 373 -1300 973 -1260
rect 2071 -740 2671 -700
rect 2071 -1260 2111 -740
rect 2631 -1260 2671 -740
rect 2071 -1300 2671 -1260
rect 3769 -740 4369 -700
rect 3769 -1260 3809 -740
rect 4329 -1260 4369 -740
rect 3769 -1300 4369 -1260
rect 5467 -740 6067 -700
rect 5467 -1260 5507 -740
rect 6027 -1260 6067 -740
rect 5467 -1300 6067 -1260
rect 7165 -740 7765 -700
rect 7165 -1260 7205 -740
rect 7725 -1260 7765 -740
rect 7165 -1300 7765 -1260
rect 8863 -740 9463 -700
rect 8863 -1260 8903 -740
rect 9423 -1260 9463 -740
rect 8863 -1300 9463 -1260
rect 10561 -740 11161 -700
rect 10561 -1260 10601 -740
rect 11121 -1260 11161 -740
rect 10561 -1300 11161 -1260
rect 12259 -740 12859 -700
rect 12259 -1260 12299 -740
rect 12819 -1260 12859 -740
rect 12259 -1300 12859 -1260
rect -13211 -1740 -12611 -1700
rect -13211 -2260 -13171 -1740
rect -12651 -2260 -12611 -1740
rect -13211 -2300 -12611 -2260
rect -11513 -1740 -10913 -1700
rect -11513 -2260 -11473 -1740
rect -10953 -2260 -10913 -1740
rect -11513 -2300 -10913 -2260
rect -9815 -1740 -9215 -1700
rect -9815 -2260 -9775 -1740
rect -9255 -2260 -9215 -1740
rect -9815 -2300 -9215 -2260
rect -8117 -1740 -7517 -1700
rect -8117 -2260 -8077 -1740
rect -7557 -2260 -7517 -1740
rect -8117 -2300 -7517 -2260
rect -6419 -1740 -5819 -1700
rect -6419 -2260 -6379 -1740
rect -5859 -2260 -5819 -1740
rect -6419 -2300 -5819 -2260
rect -4721 -1740 -4121 -1700
rect -4721 -2260 -4681 -1740
rect -4161 -2260 -4121 -1740
rect -4721 -2300 -4121 -2260
rect -3023 -1740 -2423 -1700
rect -3023 -2260 -2983 -1740
rect -2463 -2260 -2423 -1740
rect -3023 -2300 -2423 -2260
rect -1325 -1740 -725 -1700
rect -1325 -2260 -1285 -1740
rect -765 -2260 -725 -1740
rect -1325 -2300 -725 -2260
rect 373 -1740 973 -1700
rect 373 -2260 413 -1740
rect 933 -2260 973 -1740
rect 373 -2300 973 -2260
rect 2071 -1740 2671 -1700
rect 2071 -2260 2111 -1740
rect 2631 -2260 2671 -1740
rect 2071 -2300 2671 -2260
rect 3769 -1740 4369 -1700
rect 3769 -2260 3809 -1740
rect 4329 -2260 4369 -1740
rect 3769 -2300 4369 -2260
rect 5467 -1740 6067 -1700
rect 5467 -2260 5507 -1740
rect 6027 -2260 6067 -1740
rect 5467 -2300 6067 -2260
rect 7165 -1740 7765 -1700
rect 7165 -2260 7205 -1740
rect 7725 -2260 7765 -1740
rect 7165 -2300 7765 -2260
rect 8863 -1740 9463 -1700
rect 8863 -2260 8903 -1740
rect 9423 -2260 9463 -1740
rect 8863 -2300 9463 -2260
rect 10561 -1740 11161 -1700
rect 10561 -2260 10601 -1740
rect 11121 -2260 11161 -1740
rect 10561 -2300 11161 -2260
rect 12259 -1740 12859 -1700
rect 12259 -2260 12299 -1740
rect 12819 -2260 12859 -1740
rect 12259 -2300 12859 -2260
rect -13211 -2740 -12611 -2700
rect -13211 -3260 -13171 -2740
rect -12651 -3260 -12611 -2740
rect -13211 -3300 -12611 -3260
rect -11513 -2740 -10913 -2700
rect -11513 -3260 -11473 -2740
rect -10953 -3260 -10913 -2740
rect -11513 -3300 -10913 -3260
rect -9815 -2740 -9215 -2700
rect -9815 -3260 -9775 -2740
rect -9255 -3260 -9215 -2740
rect -9815 -3300 -9215 -3260
rect -8117 -2740 -7517 -2700
rect -8117 -3260 -8077 -2740
rect -7557 -3260 -7517 -2740
rect -8117 -3300 -7517 -3260
rect -6419 -2740 -5819 -2700
rect -6419 -3260 -6379 -2740
rect -5859 -3260 -5819 -2740
rect -6419 -3300 -5819 -3260
rect -4721 -2740 -4121 -2700
rect -4721 -3260 -4681 -2740
rect -4161 -3260 -4121 -2740
rect -4721 -3300 -4121 -3260
rect -3023 -2740 -2423 -2700
rect -3023 -3260 -2983 -2740
rect -2463 -3260 -2423 -2740
rect -3023 -3300 -2423 -3260
rect -1325 -2740 -725 -2700
rect -1325 -3260 -1285 -2740
rect -765 -3260 -725 -2740
rect -1325 -3300 -725 -3260
rect 373 -2740 973 -2700
rect 373 -3260 413 -2740
rect 933 -3260 973 -2740
rect 373 -3300 973 -3260
rect 2071 -2740 2671 -2700
rect 2071 -3260 2111 -2740
rect 2631 -3260 2671 -2740
rect 2071 -3300 2671 -3260
rect 3769 -2740 4369 -2700
rect 3769 -3260 3809 -2740
rect 4329 -3260 4369 -2740
rect 3769 -3300 4369 -3260
rect 5467 -2740 6067 -2700
rect 5467 -3260 5507 -2740
rect 6027 -3260 6067 -2740
rect 5467 -3300 6067 -3260
rect 7165 -2740 7765 -2700
rect 7165 -3260 7205 -2740
rect 7725 -3260 7765 -2740
rect 7165 -3300 7765 -3260
rect 8863 -2740 9463 -2700
rect 8863 -3260 8903 -2740
rect 9423 -3260 9463 -2740
rect 8863 -3300 9463 -3260
rect 10561 -2740 11161 -2700
rect 10561 -3260 10601 -2740
rect 11121 -3260 11161 -2740
rect 10561 -3300 11161 -3260
rect 12259 -2740 12859 -2700
rect 12259 -3260 12299 -2740
rect 12819 -3260 12859 -2740
rect 12259 -3300 12859 -3260
rect -13211 -3740 -12611 -3700
rect -13211 -4260 -13171 -3740
rect -12651 -4260 -12611 -3740
rect -13211 -4300 -12611 -4260
rect -11513 -3740 -10913 -3700
rect -11513 -4260 -11473 -3740
rect -10953 -4260 -10913 -3740
rect -11513 -4300 -10913 -4260
rect -9815 -3740 -9215 -3700
rect -9815 -4260 -9775 -3740
rect -9255 -4260 -9215 -3740
rect -9815 -4300 -9215 -4260
rect -8117 -3740 -7517 -3700
rect -8117 -4260 -8077 -3740
rect -7557 -4260 -7517 -3740
rect -8117 -4300 -7517 -4260
rect -6419 -3740 -5819 -3700
rect -6419 -4260 -6379 -3740
rect -5859 -4260 -5819 -3740
rect -6419 -4300 -5819 -4260
rect -4721 -3740 -4121 -3700
rect -4721 -4260 -4681 -3740
rect -4161 -4260 -4121 -3740
rect -4721 -4300 -4121 -4260
rect -3023 -3740 -2423 -3700
rect -3023 -4260 -2983 -3740
rect -2463 -4260 -2423 -3740
rect -3023 -4300 -2423 -4260
rect -1325 -3740 -725 -3700
rect -1325 -4260 -1285 -3740
rect -765 -4260 -725 -3740
rect -1325 -4300 -725 -4260
rect 373 -3740 973 -3700
rect 373 -4260 413 -3740
rect 933 -4260 973 -3740
rect 373 -4300 973 -4260
rect 2071 -3740 2671 -3700
rect 2071 -4260 2111 -3740
rect 2631 -4260 2671 -3740
rect 2071 -4300 2671 -4260
rect 3769 -3740 4369 -3700
rect 3769 -4260 3809 -3740
rect 4329 -4260 4369 -3740
rect 3769 -4300 4369 -4260
rect 5467 -3740 6067 -3700
rect 5467 -4260 5507 -3740
rect 6027 -4260 6067 -3740
rect 5467 -4300 6067 -4260
rect 7165 -3740 7765 -3700
rect 7165 -4260 7205 -3740
rect 7725 -4260 7765 -3740
rect 7165 -4300 7765 -4260
rect 8863 -3740 9463 -3700
rect 8863 -4260 8903 -3740
rect 9423 -4260 9463 -3740
rect 8863 -4300 9463 -4260
rect 10561 -3740 11161 -3700
rect 10561 -4260 10601 -3740
rect 11121 -4260 11161 -3740
rect 10561 -4300 11161 -4260
rect 12259 -3740 12859 -3700
rect 12259 -4260 12299 -3740
rect 12819 -4260 12859 -3740
rect 12259 -4300 12859 -4260
<< mimcapcontact >>
rect -13171 3740 -12651 4260
rect -11473 3740 -10953 4260
rect -9775 3740 -9255 4260
rect -8077 3740 -7557 4260
rect -6379 3740 -5859 4260
rect -4681 3740 -4161 4260
rect -2983 3740 -2463 4260
rect -1285 3740 -765 4260
rect 413 3740 933 4260
rect 2111 3740 2631 4260
rect 3809 3740 4329 4260
rect 5507 3740 6027 4260
rect 7205 3740 7725 4260
rect 8903 3740 9423 4260
rect 10601 3740 11121 4260
rect 12299 3740 12819 4260
rect -13171 2740 -12651 3260
rect -11473 2740 -10953 3260
rect -9775 2740 -9255 3260
rect -8077 2740 -7557 3260
rect -6379 2740 -5859 3260
rect -4681 2740 -4161 3260
rect -2983 2740 -2463 3260
rect -1285 2740 -765 3260
rect 413 2740 933 3260
rect 2111 2740 2631 3260
rect 3809 2740 4329 3260
rect 5507 2740 6027 3260
rect 7205 2740 7725 3260
rect 8903 2740 9423 3260
rect 10601 2740 11121 3260
rect 12299 2740 12819 3260
rect -13171 1740 -12651 2260
rect -11473 1740 -10953 2260
rect -9775 1740 -9255 2260
rect -8077 1740 -7557 2260
rect -6379 1740 -5859 2260
rect -4681 1740 -4161 2260
rect -2983 1740 -2463 2260
rect -1285 1740 -765 2260
rect 413 1740 933 2260
rect 2111 1740 2631 2260
rect 3809 1740 4329 2260
rect 5507 1740 6027 2260
rect 7205 1740 7725 2260
rect 8903 1740 9423 2260
rect 10601 1740 11121 2260
rect 12299 1740 12819 2260
rect -13171 740 -12651 1260
rect -11473 740 -10953 1260
rect -9775 740 -9255 1260
rect -8077 740 -7557 1260
rect -6379 740 -5859 1260
rect -4681 740 -4161 1260
rect -2983 740 -2463 1260
rect -1285 740 -765 1260
rect 413 740 933 1260
rect 2111 740 2631 1260
rect 3809 740 4329 1260
rect 5507 740 6027 1260
rect 7205 740 7725 1260
rect 8903 740 9423 1260
rect 10601 740 11121 1260
rect 12299 740 12819 1260
rect -13171 -260 -12651 260
rect -11473 -260 -10953 260
rect -9775 -260 -9255 260
rect -8077 -260 -7557 260
rect -6379 -260 -5859 260
rect -4681 -260 -4161 260
rect -2983 -260 -2463 260
rect -1285 -260 -765 260
rect 413 -260 933 260
rect 2111 -260 2631 260
rect 3809 -260 4329 260
rect 5507 -260 6027 260
rect 7205 -260 7725 260
rect 8903 -260 9423 260
rect 10601 -260 11121 260
rect 12299 -260 12819 260
rect -13171 -1260 -12651 -740
rect -11473 -1260 -10953 -740
rect -9775 -1260 -9255 -740
rect -8077 -1260 -7557 -740
rect -6379 -1260 -5859 -740
rect -4681 -1260 -4161 -740
rect -2983 -1260 -2463 -740
rect -1285 -1260 -765 -740
rect 413 -1260 933 -740
rect 2111 -1260 2631 -740
rect 3809 -1260 4329 -740
rect 5507 -1260 6027 -740
rect 7205 -1260 7725 -740
rect 8903 -1260 9423 -740
rect 10601 -1260 11121 -740
rect 12299 -1260 12819 -740
rect -13171 -2260 -12651 -1740
rect -11473 -2260 -10953 -1740
rect -9775 -2260 -9255 -1740
rect -8077 -2260 -7557 -1740
rect -6379 -2260 -5859 -1740
rect -4681 -2260 -4161 -1740
rect -2983 -2260 -2463 -1740
rect -1285 -2260 -765 -1740
rect 413 -2260 933 -1740
rect 2111 -2260 2631 -1740
rect 3809 -2260 4329 -1740
rect 5507 -2260 6027 -1740
rect 7205 -2260 7725 -1740
rect 8903 -2260 9423 -1740
rect 10601 -2260 11121 -1740
rect 12299 -2260 12819 -1740
rect -13171 -3260 -12651 -2740
rect -11473 -3260 -10953 -2740
rect -9775 -3260 -9255 -2740
rect -8077 -3260 -7557 -2740
rect -6379 -3260 -5859 -2740
rect -4681 -3260 -4161 -2740
rect -2983 -3260 -2463 -2740
rect -1285 -3260 -765 -2740
rect 413 -3260 933 -2740
rect 2111 -3260 2631 -2740
rect 3809 -3260 4329 -2740
rect 5507 -3260 6027 -2740
rect 7205 -3260 7725 -2740
rect 8903 -3260 9423 -2740
rect 10601 -3260 11121 -2740
rect 12299 -3260 12819 -2740
rect -13171 -4260 -12651 -3740
rect -11473 -4260 -10953 -3740
rect -9775 -4260 -9255 -3740
rect -8077 -4260 -7557 -3740
rect -6379 -4260 -5859 -3740
rect -4681 -4260 -4161 -3740
rect -2983 -4260 -2463 -3740
rect -1285 -4260 -765 -3740
rect 413 -4260 933 -3740
rect 2111 -4260 2631 -3740
rect 3809 -4260 4329 -3740
rect 5507 -4260 6027 -3740
rect 7205 -4260 7725 -3740
rect 8903 -4260 9423 -3740
rect 10601 -4260 11121 -3740
rect 12299 -4260 12819 -3740
<< metal4 >>
rect -12963 4261 -12859 4500
rect -12323 4312 -12219 4500
rect -13172 4260 -12650 4261
rect -13172 3740 -13171 4260
rect -12651 3740 -12650 4260
rect -13172 3739 -12650 3740
rect -12963 3261 -12859 3739
rect -12323 3688 -12303 4312
rect -12239 3688 -12219 4312
rect -11265 4261 -11161 4500
rect -10625 4312 -10521 4500
rect -11474 4260 -10952 4261
rect -11474 3740 -11473 4260
rect -10953 3740 -10952 4260
rect -11474 3739 -10952 3740
rect -12323 3312 -12219 3688
rect -13172 3260 -12650 3261
rect -13172 2740 -13171 3260
rect -12651 2740 -12650 3260
rect -13172 2739 -12650 2740
rect -12963 2261 -12859 2739
rect -12323 2688 -12303 3312
rect -12239 2688 -12219 3312
rect -11265 3261 -11161 3739
rect -10625 3688 -10605 4312
rect -10541 3688 -10521 4312
rect -9567 4261 -9463 4500
rect -8927 4312 -8823 4500
rect -9776 4260 -9254 4261
rect -9776 3740 -9775 4260
rect -9255 3740 -9254 4260
rect -9776 3739 -9254 3740
rect -10625 3312 -10521 3688
rect -11474 3260 -10952 3261
rect -11474 2740 -11473 3260
rect -10953 2740 -10952 3260
rect -11474 2739 -10952 2740
rect -12323 2312 -12219 2688
rect -13172 2260 -12650 2261
rect -13172 1740 -13171 2260
rect -12651 1740 -12650 2260
rect -13172 1739 -12650 1740
rect -12963 1261 -12859 1739
rect -12323 1688 -12303 2312
rect -12239 1688 -12219 2312
rect -11265 2261 -11161 2739
rect -10625 2688 -10605 3312
rect -10541 2688 -10521 3312
rect -9567 3261 -9463 3739
rect -8927 3688 -8907 4312
rect -8843 3688 -8823 4312
rect -7869 4261 -7765 4500
rect -7229 4312 -7125 4500
rect -8078 4260 -7556 4261
rect -8078 3740 -8077 4260
rect -7557 3740 -7556 4260
rect -8078 3739 -7556 3740
rect -8927 3312 -8823 3688
rect -9776 3260 -9254 3261
rect -9776 2740 -9775 3260
rect -9255 2740 -9254 3260
rect -9776 2739 -9254 2740
rect -10625 2312 -10521 2688
rect -11474 2260 -10952 2261
rect -11474 1740 -11473 2260
rect -10953 1740 -10952 2260
rect -11474 1739 -10952 1740
rect -12323 1312 -12219 1688
rect -13172 1260 -12650 1261
rect -13172 740 -13171 1260
rect -12651 740 -12650 1260
rect -13172 739 -12650 740
rect -12963 261 -12859 739
rect -12323 688 -12303 1312
rect -12239 688 -12219 1312
rect -11265 1261 -11161 1739
rect -10625 1688 -10605 2312
rect -10541 1688 -10521 2312
rect -9567 2261 -9463 2739
rect -8927 2688 -8907 3312
rect -8843 2688 -8823 3312
rect -7869 3261 -7765 3739
rect -7229 3688 -7209 4312
rect -7145 3688 -7125 4312
rect -6171 4261 -6067 4500
rect -5531 4312 -5427 4500
rect -6380 4260 -5858 4261
rect -6380 3740 -6379 4260
rect -5859 3740 -5858 4260
rect -6380 3739 -5858 3740
rect -7229 3312 -7125 3688
rect -8078 3260 -7556 3261
rect -8078 2740 -8077 3260
rect -7557 2740 -7556 3260
rect -8078 2739 -7556 2740
rect -8927 2312 -8823 2688
rect -9776 2260 -9254 2261
rect -9776 1740 -9775 2260
rect -9255 1740 -9254 2260
rect -9776 1739 -9254 1740
rect -10625 1312 -10521 1688
rect -11474 1260 -10952 1261
rect -11474 740 -11473 1260
rect -10953 740 -10952 1260
rect -11474 739 -10952 740
rect -12323 312 -12219 688
rect -13172 260 -12650 261
rect -13172 -260 -13171 260
rect -12651 -260 -12650 260
rect -13172 -261 -12650 -260
rect -12963 -739 -12859 -261
rect -12323 -312 -12303 312
rect -12239 -312 -12219 312
rect -11265 261 -11161 739
rect -10625 688 -10605 1312
rect -10541 688 -10521 1312
rect -9567 1261 -9463 1739
rect -8927 1688 -8907 2312
rect -8843 1688 -8823 2312
rect -7869 2261 -7765 2739
rect -7229 2688 -7209 3312
rect -7145 2688 -7125 3312
rect -6171 3261 -6067 3739
rect -5531 3688 -5511 4312
rect -5447 3688 -5427 4312
rect -4473 4261 -4369 4500
rect -3833 4312 -3729 4500
rect -4682 4260 -4160 4261
rect -4682 3740 -4681 4260
rect -4161 3740 -4160 4260
rect -4682 3739 -4160 3740
rect -5531 3312 -5427 3688
rect -6380 3260 -5858 3261
rect -6380 2740 -6379 3260
rect -5859 2740 -5858 3260
rect -6380 2739 -5858 2740
rect -7229 2312 -7125 2688
rect -8078 2260 -7556 2261
rect -8078 1740 -8077 2260
rect -7557 1740 -7556 2260
rect -8078 1739 -7556 1740
rect -8927 1312 -8823 1688
rect -9776 1260 -9254 1261
rect -9776 740 -9775 1260
rect -9255 740 -9254 1260
rect -9776 739 -9254 740
rect -10625 312 -10521 688
rect -11474 260 -10952 261
rect -11474 -260 -11473 260
rect -10953 -260 -10952 260
rect -11474 -261 -10952 -260
rect -12323 -688 -12219 -312
rect -13172 -740 -12650 -739
rect -13172 -1260 -13171 -740
rect -12651 -1260 -12650 -740
rect -13172 -1261 -12650 -1260
rect -12963 -1739 -12859 -1261
rect -12323 -1312 -12303 -688
rect -12239 -1312 -12219 -688
rect -11265 -739 -11161 -261
rect -10625 -312 -10605 312
rect -10541 -312 -10521 312
rect -9567 261 -9463 739
rect -8927 688 -8907 1312
rect -8843 688 -8823 1312
rect -7869 1261 -7765 1739
rect -7229 1688 -7209 2312
rect -7145 1688 -7125 2312
rect -6171 2261 -6067 2739
rect -5531 2688 -5511 3312
rect -5447 2688 -5427 3312
rect -4473 3261 -4369 3739
rect -3833 3688 -3813 4312
rect -3749 3688 -3729 4312
rect -2775 4261 -2671 4500
rect -2135 4312 -2031 4500
rect -2984 4260 -2462 4261
rect -2984 3740 -2983 4260
rect -2463 3740 -2462 4260
rect -2984 3739 -2462 3740
rect -3833 3312 -3729 3688
rect -4682 3260 -4160 3261
rect -4682 2740 -4681 3260
rect -4161 2740 -4160 3260
rect -4682 2739 -4160 2740
rect -5531 2312 -5427 2688
rect -6380 2260 -5858 2261
rect -6380 1740 -6379 2260
rect -5859 1740 -5858 2260
rect -6380 1739 -5858 1740
rect -7229 1312 -7125 1688
rect -8078 1260 -7556 1261
rect -8078 740 -8077 1260
rect -7557 740 -7556 1260
rect -8078 739 -7556 740
rect -8927 312 -8823 688
rect -9776 260 -9254 261
rect -9776 -260 -9775 260
rect -9255 -260 -9254 260
rect -9776 -261 -9254 -260
rect -10625 -688 -10521 -312
rect -11474 -740 -10952 -739
rect -11474 -1260 -11473 -740
rect -10953 -1260 -10952 -740
rect -11474 -1261 -10952 -1260
rect -12323 -1688 -12219 -1312
rect -13172 -1740 -12650 -1739
rect -13172 -2260 -13171 -1740
rect -12651 -2260 -12650 -1740
rect -13172 -2261 -12650 -2260
rect -12963 -2739 -12859 -2261
rect -12323 -2312 -12303 -1688
rect -12239 -2312 -12219 -1688
rect -11265 -1739 -11161 -1261
rect -10625 -1312 -10605 -688
rect -10541 -1312 -10521 -688
rect -9567 -739 -9463 -261
rect -8927 -312 -8907 312
rect -8843 -312 -8823 312
rect -7869 261 -7765 739
rect -7229 688 -7209 1312
rect -7145 688 -7125 1312
rect -6171 1261 -6067 1739
rect -5531 1688 -5511 2312
rect -5447 1688 -5427 2312
rect -4473 2261 -4369 2739
rect -3833 2688 -3813 3312
rect -3749 2688 -3729 3312
rect -2775 3261 -2671 3739
rect -2135 3688 -2115 4312
rect -2051 3688 -2031 4312
rect -1077 4261 -973 4500
rect -437 4312 -333 4500
rect -1286 4260 -764 4261
rect -1286 3740 -1285 4260
rect -765 3740 -764 4260
rect -1286 3739 -764 3740
rect -2135 3312 -2031 3688
rect -2984 3260 -2462 3261
rect -2984 2740 -2983 3260
rect -2463 2740 -2462 3260
rect -2984 2739 -2462 2740
rect -3833 2312 -3729 2688
rect -4682 2260 -4160 2261
rect -4682 1740 -4681 2260
rect -4161 1740 -4160 2260
rect -4682 1739 -4160 1740
rect -5531 1312 -5427 1688
rect -6380 1260 -5858 1261
rect -6380 740 -6379 1260
rect -5859 740 -5858 1260
rect -6380 739 -5858 740
rect -7229 312 -7125 688
rect -8078 260 -7556 261
rect -8078 -260 -8077 260
rect -7557 -260 -7556 260
rect -8078 -261 -7556 -260
rect -8927 -688 -8823 -312
rect -9776 -740 -9254 -739
rect -9776 -1260 -9775 -740
rect -9255 -1260 -9254 -740
rect -9776 -1261 -9254 -1260
rect -10625 -1688 -10521 -1312
rect -11474 -1740 -10952 -1739
rect -11474 -2260 -11473 -1740
rect -10953 -2260 -10952 -1740
rect -11474 -2261 -10952 -2260
rect -12323 -2688 -12219 -2312
rect -13172 -2740 -12650 -2739
rect -13172 -3260 -13171 -2740
rect -12651 -3260 -12650 -2740
rect -13172 -3261 -12650 -3260
rect -12963 -3739 -12859 -3261
rect -12323 -3312 -12303 -2688
rect -12239 -3312 -12219 -2688
rect -11265 -2739 -11161 -2261
rect -10625 -2312 -10605 -1688
rect -10541 -2312 -10521 -1688
rect -9567 -1739 -9463 -1261
rect -8927 -1312 -8907 -688
rect -8843 -1312 -8823 -688
rect -7869 -739 -7765 -261
rect -7229 -312 -7209 312
rect -7145 -312 -7125 312
rect -6171 261 -6067 739
rect -5531 688 -5511 1312
rect -5447 688 -5427 1312
rect -4473 1261 -4369 1739
rect -3833 1688 -3813 2312
rect -3749 1688 -3729 2312
rect -2775 2261 -2671 2739
rect -2135 2688 -2115 3312
rect -2051 2688 -2031 3312
rect -1077 3261 -973 3739
rect -437 3688 -417 4312
rect -353 3688 -333 4312
rect 621 4261 725 4500
rect 1261 4312 1365 4500
rect 412 4260 934 4261
rect 412 3740 413 4260
rect 933 3740 934 4260
rect 412 3739 934 3740
rect -437 3312 -333 3688
rect -1286 3260 -764 3261
rect -1286 2740 -1285 3260
rect -765 2740 -764 3260
rect -1286 2739 -764 2740
rect -2135 2312 -2031 2688
rect -2984 2260 -2462 2261
rect -2984 1740 -2983 2260
rect -2463 1740 -2462 2260
rect -2984 1739 -2462 1740
rect -3833 1312 -3729 1688
rect -4682 1260 -4160 1261
rect -4682 740 -4681 1260
rect -4161 740 -4160 1260
rect -4682 739 -4160 740
rect -5531 312 -5427 688
rect -6380 260 -5858 261
rect -6380 -260 -6379 260
rect -5859 -260 -5858 260
rect -6380 -261 -5858 -260
rect -7229 -688 -7125 -312
rect -8078 -740 -7556 -739
rect -8078 -1260 -8077 -740
rect -7557 -1260 -7556 -740
rect -8078 -1261 -7556 -1260
rect -8927 -1688 -8823 -1312
rect -9776 -1740 -9254 -1739
rect -9776 -2260 -9775 -1740
rect -9255 -2260 -9254 -1740
rect -9776 -2261 -9254 -2260
rect -10625 -2688 -10521 -2312
rect -11474 -2740 -10952 -2739
rect -11474 -3260 -11473 -2740
rect -10953 -3260 -10952 -2740
rect -11474 -3261 -10952 -3260
rect -12323 -3688 -12219 -3312
rect -13172 -3740 -12650 -3739
rect -13172 -4260 -13171 -3740
rect -12651 -4260 -12650 -3740
rect -13172 -4261 -12650 -4260
rect -12963 -4500 -12859 -4261
rect -12323 -4312 -12303 -3688
rect -12239 -4312 -12219 -3688
rect -11265 -3739 -11161 -3261
rect -10625 -3312 -10605 -2688
rect -10541 -3312 -10521 -2688
rect -9567 -2739 -9463 -2261
rect -8927 -2312 -8907 -1688
rect -8843 -2312 -8823 -1688
rect -7869 -1739 -7765 -1261
rect -7229 -1312 -7209 -688
rect -7145 -1312 -7125 -688
rect -6171 -739 -6067 -261
rect -5531 -312 -5511 312
rect -5447 -312 -5427 312
rect -4473 261 -4369 739
rect -3833 688 -3813 1312
rect -3749 688 -3729 1312
rect -2775 1261 -2671 1739
rect -2135 1688 -2115 2312
rect -2051 1688 -2031 2312
rect -1077 2261 -973 2739
rect -437 2688 -417 3312
rect -353 2688 -333 3312
rect 621 3261 725 3739
rect 1261 3688 1281 4312
rect 1345 3688 1365 4312
rect 2319 4261 2423 4500
rect 2959 4312 3063 4500
rect 2110 4260 2632 4261
rect 2110 3740 2111 4260
rect 2631 3740 2632 4260
rect 2110 3739 2632 3740
rect 1261 3312 1365 3688
rect 412 3260 934 3261
rect 412 2740 413 3260
rect 933 2740 934 3260
rect 412 2739 934 2740
rect -437 2312 -333 2688
rect -1286 2260 -764 2261
rect -1286 1740 -1285 2260
rect -765 1740 -764 2260
rect -1286 1739 -764 1740
rect -2135 1312 -2031 1688
rect -2984 1260 -2462 1261
rect -2984 740 -2983 1260
rect -2463 740 -2462 1260
rect -2984 739 -2462 740
rect -3833 312 -3729 688
rect -4682 260 -4160 261
rect -4682 -260 -4681 260
rect -4161 -260 -4160 260
rect -4682 -261 -4160 -260
rect -5531 -688 -5427 -312
rect -6380 -740 -5858 -739
rect -6380 -1260 -6379 -740
rect -5859 -1260 -5858 -740
rect -6380 -1261 -5858 -1260
rect -7229 -1688 -7125 -1312
rect -8078 -1740 -7556 -1739
rect -8078 -2260 -8077 -1740
rect -7557 -2260 -7556 -1740
rect -8078 -2261 -7556 -2260
rect -8927 -2688 -8823 -2312
rect -9776 -2740 -9254 -2739
rect -9776 -3260 -9775 -2740
rect -9255 -3260 -9254 -2740
rect -9776 -3261 -9254 -3260
rect -10625 -3688 -10521 -3312
rect -11474 -3740 -10952 -3739
rect -11474 -4260 -11473 -3740
rect -10953 -4260 -10952 -3740
rect -11474 -4261 -10952 -4260
rect -12323 -4500 -12219 -4312
rect -11265 -4500 -11161 -4261
rect -10625 -4312 -10605 -3688
rect -10541 -4312 -10521 -3688
rect -9567 -3739 -9463 -3261
rect -8927 -3312 -8907 -2688
rect -8843 -3312 -8823 -2688
rect -7869 -2739 -7765 -2261
rect -7229 -2312 -7209 -1688
rect -7145 -2312 -7125 -1688
rect -6171 -1739 -6067 -1261
rect -5531 -1312 -5511 -688
rect -5447 -1312 -5427 -688
rect -4473 -739 -4369 -261
rect -3833 -312 -3813 312
rect -3749 -312 -3729 312
rect -2775 261 -2671 739
rect -2135 688 -2115 1312
rect -2051 688 -2031 1312
rect -1077 1261 -973 1739
rect -437 1688 -417 2312
rect -353 1688 -333 2312
rect 621 2261 725 2739
rect 1261 2688 1281 3312
rect 1345 2688 1365 3312
rect 2319 3261 2423 3739
rect 2959 3688 2979 4312
rect 3043 3688 3063 4312
rect 4017 4261 4121 4500
rect 4657 4312 4761 4500
rect 3808 4260 4330 4261
rect 3808 3740 3809 4260
rect 4329 3740 4330 4260
rect 3808 3739 4330 3740
rect 2959 3312 3063 3688
rect 2110 3260 2632 3261
rect 2110 2740 2111 3260
rect 2631 2740 2632 3260
rect 2110 2739 2632 2740
rect 1261 2312 1365 2688
rect 412 2260 934 2261
rect 412 1740 413 2260
rect 933 1740 934 2260
rect 412 1739 934 1740
rect -437 1312 -333 1688
rect -1286 1260 -764 1261
rect -1286 740 -1285 1260
rect -765 740 -764 1260
rect -1286 739 -764 740
rect -2135 312 -2031 688
rect -2984 260 -2462 261
rect -2984 -260 -2983 260
rect -2463 -260 -2462 260
rect -2984 -261 -2462 -260
rect -3833 -688 -3729 -312
rect -4682 -740 -4160 -739
rect -4682 -1260 -4681 -740
rect -4161 -1260 -4160 -740
rect -4682 -1261 -4160 -1260
rect -5531 -1688 -5427 -1312
rect -6380 -1740 -5858 -1739
rect -6380 -2260 -6379 -1740
rect -5859 -2260 -5858 -1740
rect -6380 -2261 -5858 -2260
rect -7229 -2688 -7125 -2312
rect -8078 -2740 -7556 -2739
rect -8078 -3260 -8077 -2740
rect -7557 -3260 -7556 -2740
rect -8078 -3261 -7556 -3260
rect -8927 -3688 -8823 -3312
rect -9776 -3740 -9254 -3739
rect -9776 -4260 -9775 -3740
rect -9255 -4260 -9254 -3740
rect -9776 -4261 -9254 -4260
rect -10625 -4500 -10521 -4312
rect -9567 -4500 -9463 -4261
rect -8927 -4312 -8907 -3688
rect -8843 -4312 -8823 -3688
rect -7869 -3739 -7765 -3261
rect -7229 -3312 -7209 -2688
rect -7145 -3312 -7125 -2688
rect -6171 -2739 -6067 -2261
rect -5531 -2312 -5511 -1688
rect -5447 -2312 -5427 -1688
rect -4473 -1739 -4369 -1261
rect -3833 -1312 -3813 -688
rect -3749 -1312 -3729 -688
rect -2775 -739 -2671 -261
rect -2135 -312 -2115 312
rect -2051 -312 -2031 312
rect -1077 261 -973 739
rect -437 688 -417 1312
rect -353 688 -333 1312
rect 621 1261 725 1739
rect 1261 1688 1281 2312
rect 1345 1688 1365 2312
rect 2319 2261 2423 2739
rect 2959 2688 2979 3312
rect 3043 2688 3063 3312
rect 4017 3261 4121 3739
rect 4657 3688 4677 4312
rect 4741 3688 4761 4312
rect 5715 4261 5819 4500
rect 6355 4312 6459 4500
rect 5506 4260 6028 4261
rect 5506 3740 5507 4260
rect 6027 3740 6028 4260
rect 5506 3739 6028 3740
rect 4657 3312 4761 3688
rect 3808 3260 4330 3261
rect 3808 2740 3809 3260
rect 4329 2740 4330 3260
rect 3808 2739 4330 2740
rect 2959 2312 3063 2688
rect 2110 2260 2632 2261
rect 2110 1740 2111 2260
rect 2631 1740 2632 2260
rect 2110 1739 2632 1740
rect 1261 1312 1365 1688
rect 412 1260 934 1261
rect 412 740 413 1260
rect 933 740 934 1260
rect 412 739 934 740
rect -437 312 -333 688
rect -1286 260 -764 261
rect -1286 -260 -1285 260
rect -765 -260 -764 260
rect -1286 -261 -764 -260
rect -2135 -688 -2031 -312
rect -2984 -740 -2462 -739
rect -2984 -1260 -2983 -740
rect -2463 -1260 -2462 -740
rect -2984 -1261 -2462 -1260
rect -3833 -1688 -3729 -1312
rect -4682 -1740 -4160 -1739
rect -4682 -2260 -4681 -1740
rect -4161 -2260 -4160 -1740
rect -4682 -2261 -4160 -2260
rect -5531 -2688 -5427 -2312
rect -6380 -2740 -5858 -2739
rect -6380 -3260 -6379 -2740
rect -5859 -3260 -5858 -2740
rect -6380 -3261 -5858 -3260
rect -7229 -3688 -7125 -3312
rect -8078 -3740 -7556 -3739
rect -8078 -4260 -8077 -3740
rect -7557 -4260 -7556 -3740
rect -8078 -4261 -7556 -4260
rect -8927 -4500 -8823 -4312
rect -7869 -4500 -7765 -4261
rect -7229 -4312 -7209 -3688
rect -7145 -4312 -7125 -3688
rect -6171 -3739 -6067 -3261
rect -5531 -3312 -5511 -2688
rect -5447 -3312 -5427 -2688
rect -4473 -2739 -4369 -2261
rect -3833 -2312 -3813 -1688
rect -3749 -2312 -3729 -1688
rect -2775 -1739 -2671 -1261
rect -2135 -1312 -2115 -688
rect -2051 -1312 -2031 -688
rect -1077 -739 -973 -261
rect -437 -312 -417 312
rect -353 -312 -333 312
rect 621 261 725 739
rect 1261 688 1281 1312
rect 1345 688 1365 1312
rect 2319 1261 2423 1739
rect 2959 1688 2979 2312
rect 3043 1688 3063 2312
rect 4017 2261 4121 2739
rect 4657 2688 4677 3312
rect 4741 2688 4761 3312
rect 5715 3261 5819 3739
rect 6355 3688 6375 4312
rect 6439 3688 6459 4312
rect 7413 4261 7517 4500
rect 8053 4312 8157 4500
rect 7204 4260 7726 4261
rect 7204 3740 7205 4260
rect 7725 3740 7726 4260
rect 7204 3739 7726 3740
rect 6355 3312 6459 3688
rect 5506 3260 6028 3261
rect 5506 2740 5507 3260
rect 6027 2740 6028 3260
rect 5506 2739 6028 2740
rect 4657 2312 4761 2688
rect 3808 2260 4330 2261
rect 3808 1740 3809 2260
rect 4329 1740 4330 2260
rect 3808 1739 4330 1740
rect 2959 1312 3063 1688
rect 2110 1260 2632 1261
rect 2110 740 2111 1260
rect 2631 740 2632 1260
rect 2110 739 2632 740
rect 1261 312 1365 688
rect 412 260 934 261
rect 412 -260 413 260
rect 933 -260 934 260
rect 412 -261 934 -260
rect -437 -688 -333 -312
rect -1286 -740 -764 -739
rect -1286 -1260 -1285 -740
rect -765 -1260 -764 -740
rect -1286 -1261 -764 -1260
rect -2135 -1688 -2031 -1312
rect -2984 -1740 -2462 -1739
rect -2984 -2260 -2983 -1740
rect -2463 -2260 -2462 -1740
rect -2984 -2261 -2462 -2260
rect -3833 -2688 -3729 -2312
rect -4682 -2740 -4160 -2739
rect -4682 -3260 -4681 -2740
rect -4161 -3260 -4160 -2740
rect -4682 -3261 -4160 -3260
rect -5531 -3688 -5427 -3312
rect -6380 -3740 -5858 -3739
rect -6380 -4260 -6379 -3740
rect -5859 -4260 -5858 -3740
rect -6380 -4261 -5858 -4260
rect -7229 -4500 -7125 -4312
rect -6171 -4500 -6067 -4261
rect -5531 -4312 -5511 -3688
rect -5447 -4312 -5427 -3688
rect -4473 -3739 -4369 -3261
rect -3833 -3312 -3813 -2688
rect -3749 -3312 -3729 -2688
rect -2775 -2739 -2671 -2261
rect -2135 -2312 -2115 -1688
rect -2051 -2312 -2031 -1688
rect -1077 -1739 -973 -1261
rect -437 -1312 -417 -688
rect -353 -1312 -333 -688
rect 621 -739 725 -261
rect 1261 -312 1281 312
rect 1345 -312 1365 312
rect 2319 261 2423 739
rect 2959 688 2979 1312
rect 3043 688 3063 1312
rect 4017 1261 4121 1739
rect 4657 1688 4677 2312
rect 4741 1688 4761 2312
rect 5715 2261 5819 2739
rect 6355 2688 6375 3312
rect 6439 2688 6459 3312
rect 7413 3261 7517 3739
rect 8053 3688 8073 4312
rect 8137 3688 8157 4312
rect 9111 4261 9215 4500
rect 9751 4312 9855 4500
rect 8902 4260 9424 4261
rect 8902 3740 8903 4260
rect 9423 3740 9424 4260
rect 8902 3739 9424 3740
rect 8053 3312 8157 3688
rect 7204 3260 7726 3261
rect 7204 2740 7205 3260
rect 7725 2740 7726 3260
rect 7204 2739 7726 2740
rect 6355 2312 6459 2688
rect 5506 2260 6028 2261
rect 5506 1740 5507 2260
rect 6027 1740 6028 2260
rect 5506 1739 6028 1740
rect 4657 1312 4761 1688
rect 3808 1260 4330 1261
rect 3808 740 3809 1260
rect 4329 740 4330 1260
rect 3808 739 4330 740
rect 2959 312 3063 688
rect 2110 260 2632 261
rect 2110 -260 2111 260
rect 2631 -260 2632 260
rect 2110 -261 2632 -260
rect 1261 -688 1365 -312
rect 412 -740 934 -739
rect 412 -1260 413 -740
rect 933 -1260 934 -740
rect 412 -1261 934 -1260
rect -437 -1688 -333 -1312
rect -1286 -1740 -764 -1739
rect -1286 -2260 -1285 -1740
rect -765 -2260 -764 -1740
rect -1286 -2261 -764 -2260
rect -2135 -2688 -2031 -2312
rect -2984 -2740 -2462 -2739
rect -2984 -3260 -2983 -2740
rect -2463 -3260 -2462 -2740
rect -2984 -3261 -2462 -3260
rect -3833 -3688 -3729 -3312
rect -4682 -3740 -4160 -3739
rect -4682 -4260 -4681 -3740
rect -4161 -4260 -4160 -3740
rect -4682 -4261 -4160 -4260
rect -5531 -4500 -5427 -4312
rect -4473 -4500 -4369 -4261
rect -3833 -4312 -3813 -3688
rect -3749 -4312 -3729 -3688
rect -2775 -3739 -2671 -3261
rect -2135 -3312 -2115 -2688
rect -2051 -3312 -2031 -2688
rect -1077 -2739 -973 -2261
rect -437 -2312 -417 -1688
rect -353 -2312 -333 -1688
rect 621 -1739 725 -1261
rect 1261 -1312 1281 -688
rect 1345 -1312 1365 -688
rect 2319 -739 2423 -261
rect 2959 -312 2979 312
rect 3043 -312 3063 312
rect 4017 261 4121 739
rect 4657 688 4677 1312
rect 4741 688 4761 1312
rect 5715 1261 5819 1739
rect 6355 1688 6375 2312
rect 6439 1688 6459 2312
rect 7413 2261 7517 2739
rect 8053 2688 8073 3312
rect 8137 2688 8157 3312
rect 9111 3261 9215 3739
rect 9751 3688 9771 4312
rect 9835 3688 9855 4312
rect 10809 4261 10913 4500
rect 11449 4312 11553 4500
rect 10600 4260 11122 4261
rect 10600 3740 10601 4260
rect 11121 3740 11122 4260
rect 10600 3739 11122 3740
rect 9751 3312 9855 3688
rect 8902 3260 9424 3261
rect 8902 2740 8903 3260
rect 9423 2740 9424 3260
rect 8902 2739 9424 2740
rect 8053 2312 8157 2688
rect 7204 2260 7726 2261
rect 7204 1740 7205 2260
rect 7725 1740 7726 2260
rect 7204 1739 7726 1740
rect 6355 1312 6459 1688
rect 5506 1260 6028 1261
rect 5506 740 5507 1260
rect 6027 740 6028 1260
rect 5506 739 6028 740
rect 4657 312 4761 688
rect 3808 260 4330 261
rect 3808 -260 3809 260
rect 4329 -260 4330 260
rect 3808 -261 4330 -260
rect 2959 -688 3063 -312
rect 2110 -740 2632 -739
rect 2110 -1260 2111 -740
rect 2631 -1260 2632 -740
rect 2110 -1261 2632 -1260
rect 1261 -1688 1365 -1312
rect 412 -1740 934 -1739
rect 412 -2260 413 -1740
rect 933 -2260 934 -1740
rect 412 -2261 934 -2260
rect -437 -2688 -333 -2312
rect -1286 -2740 -764 -2739
rect -1286 -3260 -1285 -2740
rect -765 -3260 -764 -2740
rect -1286 -3261 -764 -3260
rect -2135 -3688 -2031 -3312
rect -2984 -3740 -2462 -3739
rect -2984 -4260 -2983 -3740
rect -2463 -4260 -2462 -3740
rect -2984 -4261 -2462 -4260
rect -3833 -4500 -3729 -4312
rect -2775 -4500 -2671 -4261
rect -2135 -4312 -2115 -3688
rect -2051 -4312 -2031 -3688
rect -1077 -3739 -973 -3261
rect -437 -3312 -417 -2688
rect -353 -3312 -333 -2688
rect 621 -2739 725 -2261
rect 1261 -2312 1281 -1688
rect 1345 -2312 1365 -1688
rect 2319 -1739 2423 -1261
rect 2959 -1312 2979 -688
rect 3043 -1312 3063 -688
rect 4017 -739 4121 -261
rect 4657 -312 4677 312
rect 4741 -312 4761 312
rect 5715 261 5819 739
rect 6355 688 6375 1312
rect 6439 688 6459 1312
rect 7413 1261 7517 1739
rect 8053 1688 8073 2312
rect 8137 1688 8157 2312
rect 9111 2261 9215 2739
rect 9751 2688 9771 3312
rect 9835 2688 9855 3312
rect 10809 3261 10913 3739
rect 11449 3688 11469 4312
rect 11533 3688 11553 4312
rect 12507 4261 12611 4500
rect 13147 4312 13251 4500
rect 12298 4260 12820 4261
rect 12298 3740 12299 4260
rect 12819 3740 12820 4260
rect 12298 3739 12820 3740
rect 11449 3312 11553 3688
rect 10600 3260 11122 3261
rect 10600 2740 10601 3260
rect 11121 2740 11122 3260
rect 10600 2739 11122 2740
rect 9751 2312 9855 2688
rect 8902 2260 9424 2261
rect 8902 1740 8903 2260
rect 9423 1740 9424 2260
rect 8902 1739 9424 1740
rect 8053 1312 8157 1688
rect 7204 1260 7726 1261
rect 7204 740 7205 1260
rect 7725 740 7726 1260
rect 7204 739 7726 740
rect 6355 312 6459 688
rect 5506 260 6028 261
rect 5506 -260 5507 260
rect 6027 -260 6028 260
rect 5506 -261 6028 -260
rect 4657 -688 4761 -312
rect 3808 -740 4330 -739
rect 3808 -1260 3809 -740
rect 4329 -1260 4330 -740
rect 3808 -1261 4330 -1260
rect 2959 -1688 3063 -1312
rect 2110 -1740 2632 -1739
rect 2110 -2260 2111 -1740
rect 2631 -2260 2632 -1740
rect 2110 -2261 2632 -2260
rect 1261 -2688 1365 -2312
rect 412 -2740 934 -2739
rect 412 -3260 413 -2740
rect 933 -3260 934 -2740
rect 412 -3261 934 -3260
rect -437 -3688 -333 -3312
rect -1286 -3740 -764 -3739
rect -1286 -4260 -1285 -3740
rect -765 -4260 -764 -3740
rect -1286 -4261 -764 -4260
rect -2135 -4500 -2031 -4312
rect -1077 -4500 -973 -4261
rect -437 -4312 -417 -3688
rect -353 -4312 -333 -3688
rect 621 -3739 725 -3261
rect 1261 -3312 1281 -2688
rect 1345 -3312 1365 -2688
rect 2319 -2739 2423 -2261
rect 2959 -2312 2979 -1688
rect 3043 -2312 3063 -1688
rect 4017 -1739 4121 -1261
rect 4657 -1312 4677 -688
rect 4741 -1312 4761 -688
rect 5715 -739 5819 -261
rect 6355 -312 6375 312
rect 6439 -312 6459 312
rect 7413 261 7517 739
rect 8053 688 8073 1312
rect 8137 688 8157 1312
rect 9111 1261 9215 1739
rect 9751 1688 9771 2312
rect 9835 1688 9855 2312
rect 10809 2261 10913 2739
rect 11449 2688 11469 3312
rect 11533 2688 11553 3312
rect 12507 3261 12611 3739
rect 13147 3688 13167 4312
rect 13231 3688 13251 4312
rect 13147 3312 13251 3688
rect 12298 3260 12820 3261
rect 12298 2740 12299 3260
rect 12819 2740 12820 3260
rect 12298 2739 12820 2740
rect 11449 2312 11553 2688
rect 10600 2260 11122 2261
rect 10600 1740 10601 2260
rect 11121 1740 11122 2260
rect 10600 1739 11122 1740
rect 9751 1312 9855 1688
rect 8902 1260 9424 1261
rect 8902 740 8903 1260
rect 9423 740 9424 1260
rect 8902 739 9424 740
rect 8053 312 8157 688
rect 7204 260 7726 261
rect 7204 -260 7205 260
rect 7725 -260 7726 260
rect 7204 -261 7726 -260
rect 6355 -688 6459 -312
rect 5506 -740 6028 -739
rect 5506 -1260 5507 -740
rect 6027 -1260 6028 -740
rect 5506 -1261 6028 -1260
rect 4657 -1688 4761 -1312
rect 3808 -1740 4330 -1739
rect 3808 -2260 3809 -1740
rect 4329 -2260 4330 -1740
rect 3808 -2261 4330 -2260
rect 2959 -2688 3063 -2312
rect 2110 -2740 2632 -2739
rect 2110 -3260 2111 -2740
rect 2631 -3260 2632 -2740
rect 2110 -3261 2632 -3260
rect 1261 -3688 1365 -3312
rect 412 -3740 934 -3739
rect 412 -4260 413 -3740
rect 933 -4260 934 -3740
rect 412 -4261 934 -4260
rect -437 -4500 -333 -4312
rect 621 -4500 725 -4261
rect 1261 -4312 1281 -3688
rect 1345 -4312 1365 -3688
rect 2319 -3739 2423 -3261
rect 2959 -3312 2979 -2688
rect 3043 -3312 3063 -2688
rect 4017 -2739 4121 -2261
rect 4657 -2312 4677 -1688
rect 4741 -2312 4761 -1688
rect 5715 -1739 5819 -1261
rect 6355 -1312 6375 -688
rect 6439 -1312 6459 -688
rect 7413 -739 7517 -261
rect 8053 -312 8073 312
rect 8137 -312 8157 312
rect 9111 261 9215 739
rect 9751 688 9771 1312
rect 9835 688 9855 1312
rect 10809 1261 10913 1739
rect 11449 1688 11469 2312
rect 11533 1688 11553 2312
rect 12507 2261 12611 2739
rect 13147 2688 13167 3312
rect 13231 2688 13251 3312
rect 13147 2312 13251 2688
rect 12298 2260 12820 2261
rect 12298 1740 12299 2260
rect 12819 1740 12820 2260
rect 12298 1739 12820 1740
rect 11449 1312 11553 1688
rect 10600 1260 11122 1261
rect 10600 740 10601 1260
rect 11121 740 11122 1260
rect 10600 739 11122 740
rect 9751 312 9855 688
rect 8902 260 9424 261
rect 8902 -260 8903 260
rect 9423 -260 9424 260
rect 8902 -261 9424 -260
rect 8053 -688 8157 -312
rect 7204 -740 7726 -739
rect 7204 -1260 7205 -740
rect 7725 -1260 7726 -740
rect 7204 -1261 7726 -1260
rect 6355 -1688 6459 -1312
rect 5506 -1740 6028 -1739
rect 5506 -2260 5507 -1740
rect 6027 -2260 6028 -1740
rect 5506 -2261 6028 -2260
rect 4657 -2688 4761 -2312
rect 3808 -2740 4330 -2739
rect 3808 -3260 3809 -2740
rect 4329 -3260 4330 -2740
rect 3808 -3261 4330 -3260
rect 2959 -3688 3063 -3312
rect 2110 -3740 2632 -3739
rect 2110 -4260 2111 -3740
rect 2631 -4260 2632 -3740
rect 2110 -4261 2632 -4260
rect 1261 -4500 1365 -4312
rect 2319 -4500 2423 -4261
rect 2959 -4312 2979 -3688
rect 3043 -4312 3063 -3688
rect 4017 -3739 4121 -3261
rect 4657 -3312 4677 -2688
rect 4741 -3312 4761 -2688
rect 5715 -2739 5819 -2261
rect 6355 -2312 6375 -1688
rect 6439 -2312 6459 -1688
rect 7413 -1739 7517 -1261
rect 8053 -1312 8073 -688
rect 8137 -1312 8157 -688
rect 9111 -739 9215 -261
rect 9751 -312 9771 312
rect 9835 -312 9855 312
rect 10809 261 10913 739
rect 11449 688 11469 1312
rect 11533 688 11553 1312
rect 12507 1261 12611 1739
rect 13147 1688 13167 2312
rect 13231 1688 13251 2312
rect 13147 1312 13251 1688
rect 12298 1260 12820 1261
rect 12298 740 12299 1260
rect 12819 740 12820 1260
rect 12298 739 12820 740
rect 11449 312 11553 688
rect 10600 260 11122 261
rect 10600 -260 10601 260
rect 11121 -260 11122 260
rect 10600 -261 11122 -260
rect 9751 -688 9855 -312
rect 8902 -740 9424 -739
rect 8902 -1260 8903 -740
rect 9423 -1260 9424 -740
rect 8902 -1261 9424 -1260
rect 8053 -1688 8157 -1312
rect 7204 -1740 7726 -1739
rect 7204 -2260 7205 -1740
rect 7725 -2260 7726 -1740
rect 7204 -2261 7726 -2260
rect 6355 -2688 6459 -2312
rect 5506 -2740 6028 -2739
rect 5506 -3260 5507 -2740
rect 6027 -3260 6028 -2740
rect 5506 -3261 6028 -3260
rect 4657 -3688 4761 -3312
rect 3808 -3740 4330 -3739
rect 3808 -4260 3809 -3740
rect 4329 -4260 4330 -3740
rect 3808 -4261 4330 -4260
rect 2959 -4500 3063 -4312
rect 4017 -4500 4121 -4261
rect 4657 -4312 4677 -3688
rect 4741 -4312 4761 -3688
rect 5715 -3739 5819 -3261
rect 6355 -3312 6375 -2688
rect 6439 -3312 6459 -2688
rect 7413 -2739 7517 -2261
rect 8053 -2312 8073 -1688
rect 8137 -2312 8157 -1688
rect 9111 -1739 9215 -1261
rect 9751 -1312 9771 -688
rect 9835 -1312 9855 -688
rect 10809 -739 10913 -261
rect 11449 -312 11469 312
rect 11533 -312 11553 312
rect 12507 261 12611 739
rect 13147 688 13167 1312
rect 13231 688 13251 1312
rect 13147 312 13251 688
rect 12298 260 12820 261
rect 12298 -260 12299 260
rect 12819 -260 12820 260
rect 12298 -261 12820 -260
rect 11449 -688 11553 -312
rect 10600 -740 11122 -739
rect 10600 -1260 10601 -740
rect 11121 -1260 11122 -740
rect 10600 -1261 11122 -1260
rect 9751 -1688 9855 -1312
rect 8902 -1740 9424 -1739
rect 8902 -2260 8903 -1740
rect 9423 -2260 9424 -1740
rect 8902 -2261 9424 -2260
rect 8053 -2688 8157 -2312
rect 7204 -2740 7726 -2739
rect 7204 -3260 7205 -2740
rect 7725 -3260 7726 -2740
rect 7204 -3261 7726 -3260
rect 6355 -3688 6459 -3312
rect 5506 -3740 6028 -3739
rect 5506 -4260 5507 -3740
rect 6027 -4260 6028 -3740
rect 5506 -4261 6028 -4260
rect 4657 -4500 4761 -4312
rect 5715 -4500 5819 -4261
rect 6355 -4312 6375 -3688
rect 6439 -4312 6459 -3688
rect 7413 -3739 7517 -3261
rect 8053 -3312 8073 -2688
rect 8137 -3312 8157 -2688
rect 9111 -2739 9215 -2261
rect 9751 -2312 9771 -1688
rect 9835 -2312 9855 -1688
rect 10809 -1739 10913 -1261
rect 11449 -1312 11469 -688
rect 11533 -1312 11553 -688
rect 12507 -739 12611 -261
rect 13147 -312 13167 312
rect 13231 -312 13251 312
rect 13147 -688 13251 -312
rect 12298 -740 12820 -739
rect 12298 -1260 12299 -740
rect 12819 -1260 12820 -740
rect 12298 -1261 12820 -1260
rect 11449 -1688 11553 -1312
rect 10600 -1740 11122 -1739
rect 10600 -2260 10601 -1740
rect 11121 -2260 11122 -1740
rect 10600 -2261 11122 -2260
rect 9751 -2688 9855 -2312
rect 8902 -2740 9424 -2739
rect 8902 -3260 8903 -2740
rect 9423 -3260 9424 -2740
rect 8902 -3261 9424 -3260
rect 8053 -3688 8157 -3312
rect 7204 -3740 7726 -3739
rect 7204 -4260 7205 -3740
rect 7725 -4260 7726 -3740
rect 7204 -4261 7726 -4260
rect 6355 -4500 6459 -4312
rect 7413 -4500 7517 -4261
rect 8053 -4312 8073 -3688
rect 8137 -4312 8157 -3688
rect 9111 -3739 9215 -3261
rect 9751 -3312 9771 -2688
rect 9835 -3312 9855 -2688
rect 10809 -2739 10913 -2261
rect 11449 -2312 11469 -1688
rect 11533 -2312 11553 -1688
rect 12507 -1739 12611 -1261
rect 13147 -1312 13167 -688
rect 13231 -1312 13251 -688
rect 13147 -1688 13251 -1312
rect 12298 -1740 12820 -1739
rect 12298 -2260 12299 -1740
rect 12819 -2260 12820 -1740
rect 12298 -2261 12820 -2260
rect 11449 -2688 11553 -2312
rect 10600 -2740 11122 -2739
rect 10600 -3260 10601 -2740
rect 11121 -3260 11122 -2740
rect 10600 -3261 11122 -3260
rect 9751 -3688 9855 -3312
rect 8902 -3740 9424 -3739
rect 8902 -4260 8903 -3740
rect 9423 -4260 9424 -3740
rect 8902 -4261 9424 -4260
rect 8053 -4500 8157 -4312
rect 9111 -4500 9215 -4261
rect 9751 -4312 9771 -3688
rect 9835 -4312 9855 -3688
rect 10809 -3739 10913 -3261
rect 11449 -3312 11469 -2688
rect 11533 -3312 11553 -2688
rect 12507 -2739 12611 -2261
rect 13147 -2312 13167 -1688
rect 13231 -2312 13251 -1688
rect 13147 -2688 13251 -2312
rect 12298 -2740 12820 -2739
rect 12298 -3260 12299 -2740
rect 12819 -3260 12820 -2740
rect 12298 -3261 12820 -3260
rect 11449 -3688 11553 -3312
rect 10600 -3740 11122 -3739
rect 10600 -4260 10601 -3740
rect 11121 -4260 11122 -3740
rect 10600 -4261 11122 -4260
rect 9751 -4500 9855 -4312
rect 10809 -4500 10913 -4261
rect 11449 -4312 11469 -3688
rect 11533 -4312 11553 -3688
rect 12507 -3739 12611 -3261
rect 13147 -3312 13167 -2688
rect 13231 -3312 13251 -2688
rect 13147 -3688 13251 -3312
rect 12298 -3740 12820 -3739
rect 12298 -4260 12299 -3740
rect 12819 -4260 12820 -3740
rect 12298 -4261 12820 -4260
rect 11449 -4500 11553 -4312
rect 12507 -4500 12611 -4261
rect 13147 -4312 13167 -3688
rect 13231 -4312 13251 -3688
rect 13147 -4500 13251 -4312
<< labels >>
rlabel via3 -12271 -4000 -12271 -4000 0 C2_0
port 1 nsew
rlabel mimcapcontact -12911 -4000 -12911 -4000 0 C1_0
port 2 nsew
rlabel via3 -10573 -4000 -10573 -4000 0 C2_1
port 3 nsew
rlabel mimcapcontact -11213 -4000 -11213 -4000 0 C1_1
port 4 nsew
rlabel via3 -8875 -4000 -8875 -4000 0 C2_2
port 5 nsew
rlabel mimcapcontact -9515 -4000 -9515 -4000 0 C1_2
port 6 nsew
rlabel via3 -7177 -4000 -7177 -4000 0 C2_3
port 7 nsew
rlabel mimcapcontact -7817 -4000 -7817 -4000 0 C1_3
port 8 nsew
rlabel via3 -5479 -4000 -5479 -4000 0 C2_4
port 9 nsew
rlabel mimcapcontact -6119 -4000 -6119 -4000 0 C1_4
port 10 nsew
rlabel via3 -3781 -4000 -3781 -4000 0 C2_5
port 11 nsew
rlabel mimcapcontact -4421 -4000 -4421 -4000 0 C1_5
port 12 nsew
rlabel via3 -2083 -4000 -2083 -4000 0 C2_6
port 13 nsew
rlabel mimcapcontact -2723 -4000 -2723 -4000 0 C1_6
port 14 nsew
rlabel via3 -385 -4000 -385 -4000 0 C2_7
port 15 nsew
rlabel mimcapcontact -1025 -4000 -1025 -4000 0 C1_7
port 16 nsew
rlabel via3 1313 -4000 1313 -4000 0 C2_8
port 17 nsew
rlabel mimcapcontact 673 -4000 673 -4000 0 C1_8
port 18 nsew
rlabel via3 3011 -4000 3011 -4000 0 C2_9
port 19 nsew
rlabel mimcapcontact 2371 -4000 2371 -4000 0 C1_9
port 20 nsew
rlabel via3 4709 -4000 4709 -4000 0 C2_10
port 21 nsew
rlabel mimcapcontact 4069 -4000 4069 -4000 0 C1_10
port 22 nsew
rlabel via3 6407 -4000 6407 -4000 0 C2_11
port 23 nsew
rlabel mimcapcontact 5767 -4000 5767 -4000 0 C1_11
port 24 nsew
rlabel via3 8105 -4000 8105 -4000 0 C2_12
port 25 nsew
rlabel mimcapcontact 7465 -4000 7465 -4000 0 C1_12
port 26 nsew
rlabel via3 9803 -4000 9803 -4000 0 C2_13
port 27 nsew
rlabel mimcapcontact 9163 -4000 9163 -4000 0 C1_13
port 28 nsew
rlabel via3 11501 -4000 11501 -4000 0 C2_14
port 29 nsew
rlabel mimcapcontact 10861 -4000 10861 -4000 0 C1_14
port 30 nsew
rlabel via3 13199 -4000 13199 -4000 0 C2_15
port 31 nsew
rlabel mimcapcontact 12559 -4000 12559 -4000 0 C1_15
port 32 nsew
<< properties >>
string FIXED_BBOX 12219 3660 12899 4340
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 3 l 3 val 20.28 carea 2.00 cperi 0.19 class capacitor nx 16 ny 9 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100 stack 1 doports 1
<< end >>
