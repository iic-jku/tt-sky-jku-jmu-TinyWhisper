* PEX produced on Sun Nov  9 08:18:58 PM CET 2025 using /foss/tools/sak/iic-pex.sh with m=1 and s=1
* NGSPICE file created from iq_modulator.ext - technology: sky130A

.subckt iq_modulator_pex vout_RF vinn_I vinp_I vinp_Q vinn_Q VSS VDD di_LO_IX di_LO_I
+ di_LO_QX di_LO_Q di_afe_en
X0 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout C3_1x5_3.bottom VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl C3_1x5_1.bottom VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2 VSS iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3 VSS di_afe_en iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X4 di_LO_I VDD iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X5 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout C3_1x5_1.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X6 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_123 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_124 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X7 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X8 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X9 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X10 VDD iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X11 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X12 VSS iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X13 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X14 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_80 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_79 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X15 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X16 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 C3_1x5_1.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X17 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X18 VSS iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X19 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=279.66 ps=1.9598k w=3 l=0.15
X20 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X21 C2_3x7_2.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_37 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X22 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_112 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_111 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X23 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=18.4 ps=148.8 w=1 l=0.15
X24 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n C3_1x5_3.bottom VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X25 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_26 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_27 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X26 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X27 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X28 C3_1x5_1.bottom C3_1x5_1.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X29 C3_1x5_1.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X30 C2_3x7_2.top C2_3x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X31 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_113 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_114 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X32 C3_1x5_1.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl C3_1x5_1.bottom VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=29.46 ps=204.67999 w=3 l=0.15
X33 VDD iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=3.81 ps=8.54 w=3 l=0.15
X34 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_75 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_74 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X35 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X36 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X37 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X38 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_29 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_28 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X39 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X40 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl C3_1x5_3.bottom VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X41 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_101 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_102 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X42 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_53 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_52 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X43 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_87 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_88 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X44 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X45 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X46 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_73 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_74 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X47 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_39 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_38 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X48 VDD iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X49 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X50 C3_1x5_1.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl C3_1x5_1.bottom VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X51 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_127 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_128 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X52 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_127 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_126 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X53 iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X54 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 C3_1x5_3.top C3_1x5_3.bottom VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X55 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X56 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X57 C3_1x5_1.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X58 C2_3x7_2.top C2_3x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X59 C3_1x5_1.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n C3_1x5_1.bottom VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=9.82 ps=76.68 w=1 l=0.15
X60 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X61 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X62 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VSS di_LO_QX VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.93 ps=6.62 w=3 l=0.15
X63 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X64 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout C3_1x5_3.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X65 iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X66 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X67 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_112 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_113 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X68 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X69 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_109 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_110 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X70 C3_1x5_1.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n C3_1x5_1.bottom VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X71 VDD iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X72 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_102 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_103 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X73 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X74 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X75 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_25 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_24 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X76 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X77 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=55.2 ps=372.79999 w=3 l=0.15
X78 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X79 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X80 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X81 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=0 ps=0 w=9 l=1
X82 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_11 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_12 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X83 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X84 VSS iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X85 VSS iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X86 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=93.22 ps=735.79999 w=1 l=0.15
X87 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X88 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_50 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_49 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X89 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n C3_1x5_1.bottom VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X90 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_91 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_92 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X91 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_11 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_10 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X92 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X93 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X94 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_72 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_71 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X95 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_105 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_104 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X96 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_91 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_90 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X97 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X98 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X99 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X100 VDD iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X101 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_35 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X102 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_70 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_71 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X103 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X104 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_124 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_125 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X105 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X106 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl C3_1x5_1.bottom VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X107 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X108 iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X109 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X110 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X111 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_124 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_123 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X112 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X113 VDD di_LO_IX iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X114 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VDD di_LO_QX VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X115 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X116 C3_1x5_1.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X117 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X118 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_132 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_133 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X119 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X120 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X121 C2_3x7_2.top C2_3x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X122 iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X123 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin di_LO_IX VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X124 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X125 VSS iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X126 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X127 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_15 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_14 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X128 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VSS di_LO_I VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.93 ps=6.62 w=3 l=0.15
X129 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X130 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_0 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X131 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X132 C3_1x5_1.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X133 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X134 C3_1x5_3.bottom C3_1x5_3.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X135 VSS VDD iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X136 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=29.46 ps=204.67999 w=3 l=0.15
X137 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_75 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_76 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X138 iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X139 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X140 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_13 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_14 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X141 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_117 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_116 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X142 VDD iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X143 iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X144 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_30 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_31 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X145 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_74 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_75 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X146 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X147 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_107 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_108 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X148 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_65 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_66 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X149 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X150 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X151 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_102 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_101 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X152 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X153 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_58 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_59 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X154 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_52 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_53 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X155 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_38 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_39 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X156 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_88 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_87 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X157 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=0 ps=0 w=9 l=1
X158 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X159 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_74 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_73 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X160 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X161 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X162 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_23 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_22 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X163 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_128 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_127 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X164 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X165 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X166 C3_1x5_1.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X167 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X168 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X169 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X170 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n di_afe_en VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X171 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=0 ps=0 w=9 l=1
X172 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X173 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_6 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_5 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X174 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X175 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X176 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X177 C3_1x5_1.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X178 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X179 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X180 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X181 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=9.82 ps=76.68 w=1 l=0.15
X182 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_31 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_32 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X183 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_96 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_97 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X184 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X185 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_67 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_66 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X186 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X187 VSS iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X188 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X189 VSS iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X190 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X191 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_12 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_11 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X192 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n di_afe_en VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X193 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X194 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X195 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X196 VDD iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X197 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X198 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_92 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_91 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X199 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_10 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_11 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X200 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_98 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X201 VDD iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X202 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X203 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X204 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout C3_1x5_3.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X205 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_104 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_105 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X206 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_90 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_91 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X207 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X208 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_13 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_14 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X209 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_89 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_88 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X210 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X211 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n C3_1x5_1.bottom VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X212 VSS VDD iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X213 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X214 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X215 C3_1x5_3.bottom C3_1x5_3.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X216 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_45 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_46 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X217 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_3 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_4 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X218 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X219 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X220 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X221 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_114 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_113 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X222 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X223 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X224 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X225 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X226 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_35 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X227 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X228 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X229 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl C3_1x5_1.bottom VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X230 C2_3x7_2.bottom C2_3x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X231 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_28 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_29 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X232 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X233 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X234 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_126 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_127 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X235 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X236 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X237 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X238 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=29.46 ps=204.67999 w=3 l=0.15
X239 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X240 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_14 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_15 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X241 VSS iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=1.27 ps=4.54 w=1 l=0.15
X242 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_0 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_1 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X243 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout C3_1x5_1.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X244 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X245 iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X246 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X247 C3_1x5_1.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X248 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_14 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_13 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X249 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_110 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_109 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X250 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_129 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_128 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X251 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_116 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_117 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X252 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X253 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X254 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_69 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_70 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X255 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X256 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 C3_1x5_3.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X257 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X258 C3_1x5_3.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X259 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X260 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X261 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_24 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_25 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X262 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X263 iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X264 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_119 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_118 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X265 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X266 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_101 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_102 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X267 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_59 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_60 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X268 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X269 VSS iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=1.27 ps=4.54 w=1 l=0.15
X270 VSS VDD iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X271 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_16 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X272 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X273 di_LO_IX VDD iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X274 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X275 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X276 C3_1x5_3.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X277 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X278 VDD iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X279 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_77 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_78 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X280 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X281 C3_1x5_1.top C3_1x5_1.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X282 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X283 VSS VDD iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X284 VSS iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X285 C2_3x7_2.bottom C2_3x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X286 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_131 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_130 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X287 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_32 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_31 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X288 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_66 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_67 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X289 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X290 iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X291 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n C3_1x5_1.bottom VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X292 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X293 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_61 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_60 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X294 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X295 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X296 VDD iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=3.81 ps=8.54 w=3 l=0.15
X297 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X298 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X299 VSS iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=1.27 ps=4.54 w=1 l=0.15
X300 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_93 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_92 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X301 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 C3_1x5_1.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X302 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl C3_1x5_1.bottom VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X303 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_131 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_132 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X304 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X305 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout C3_1x5_1.bottom VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X306 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X307 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_7 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_8 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X308 VDD iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X309 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_83 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_82 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X310 C2_3x7_2.bottom C2_3x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X311 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VSS di_LO_Q VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.93 ps=6.62 w=3 l=0.15
X312 VSS VDD iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X313 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X314 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_76 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_75 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X315 C2_3x7_2.bottom C2_3x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X316 VSS iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X317 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_95 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_94 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X318 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_39 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_40 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X319 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_81 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_80 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X320 C2_3x7_2.top C2_3x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X321 VDD iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X322 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_66 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_65 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X323 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X324 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_108 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_107 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X325 iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X326 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_107 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_108 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X327 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X328 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_93 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_94 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X329 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_29 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_30 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X330 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_133 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_134 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X331 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_22 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_23 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X332 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin di_LO_QX VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X333 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X334 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X335 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X336 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X337 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X338 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X339 C2_3x7_2.top C2_3x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X340 C3_1x5_3.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X341 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X342 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X343 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X344 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X345 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X346 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_123 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_122 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X347 C3_1x5_3.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl C3_1x5_3.bottom VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=29.46 ps=204.67999 w=3 l=0.15
X348 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X349 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X350 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 C3_1x5_1.top C3_1x5_1.bottom VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X351 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_73 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_74 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X352 C1_5x7_2.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_18 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X353 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_3 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_4 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X354 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X355 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X356 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X357 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_111 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_112 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X358 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_105 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_106 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X359 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_97 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_98 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X360 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_119 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_120 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X361 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout C3_1x5_1.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X362 C3_1x5_3.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n C3_1x5_3.bottom VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=9.82 ps=76.68 w=1 l=0.15
X363 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 C3_1x5_1.top C3_1x5_1.bottom VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X364 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_98 C3_1x5_3.top VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X365 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_78 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_77 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X366 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X367 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VDD di_LO_Q VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X368 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_111 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_110 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X369 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 C3_1x5_3.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X370 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_21 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_20 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X371 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X372 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X373 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X374 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X375 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X376 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_14 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_13 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X377 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_88 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_89 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X378 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X379 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X380 VDD iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=3.81 ps=8.54 w=3 l=0.15
X381 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X382 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X383 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_53 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_52 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X384 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_130 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_131 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X385 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X386 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout C3_1x5_1.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X387 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X388 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_4 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_3 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X389 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VSS di_LO_IX VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.93 ps=6.62 w=3 l=0.15
X390 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_46 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_45 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X391 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X392 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X393 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X394 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X395 C2_3x7_2.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_35 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X396 iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X397 VDD iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X398 iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X399 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_57 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_56 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X400 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_21 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_22 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X401 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_55 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_54 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X402 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=9.82 ps=76.68 w=1 l=0.15
X403 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X404 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout C3_1x5_3.bottom VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X405 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X406 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X407 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_35 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_34 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X408 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_69 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_70 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X409 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_21 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_20 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X410 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_55 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_56 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X411 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X412 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_87 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_86 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X413 C2_3x7_2.top C2_3x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X414 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X415 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X416 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X417 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X418 C3_1x5_3.top C3_1x5_3.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X419 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_135 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_136 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X420 C3_1x5_1.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_136 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X421 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_2 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X422 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_123 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_122 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X423 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_77 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_76 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X424 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X425 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_128 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_129 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X426 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_94 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_95 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X427 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_80 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_81 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X428 C3_1x5_1.bottom C3_1x5_1.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X429 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_70 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_69 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X430 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X431 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X432 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X433 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X434 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X435 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_118 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_119 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X436 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_108 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_107 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X437 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_94 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_93 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X438 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_43 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_44 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X439 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X440 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X441 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_102 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_101 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X442 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_60 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_59 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X443 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_134 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_133 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X444 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X445 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X446 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X447 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_16 C1_5x7_2.top VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X448 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_33 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_34 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X449 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X450 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X451 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X452 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X453 VDD iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X454 VSS VDD iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X455 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X456 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X457 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X458 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X459 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X460 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_25 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_24 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X461 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X462 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_51 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_52 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X463 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_87 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_86 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X464 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_37 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_38 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X465 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X466 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_73 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_72 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X467 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_127 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_126 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X468 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_117 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_116 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X469 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout C3_1x5_1.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X470 VDD iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X471 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_18 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X472 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X473 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_4 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_3 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X474 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X475 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X476 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_67 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_68 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X477 C2_3x7_2.top C2_3x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X478 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout C3_1x5_3.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X479 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n C3_1x5_3.bottom VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X480 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 C3_1x5_3.top C3_1x5_3.bottom VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X481 VDD iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X482 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X483 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_112 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_111 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X484 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_98 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_97 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X485 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_60 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_61 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X486 VSS iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=1.27 ps=4.54 w=1 l=0.15
X487 VDD iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X488 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_120 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_119 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X489 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X490 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X491 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X492 iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X493 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_100 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X494 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X495 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X496 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_110 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_111 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X497 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X498 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_92 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_93 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X499 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_132 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_131 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X500 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X501 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_15 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_14 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X502 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X503 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout C3_1x5_3.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X504 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X505 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl C3_1x5_3.bottom VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X506 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_8 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_7 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X507 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X508 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_82 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_83 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X509 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X510 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X511 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X512 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X513 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout C3_1x5_1.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X514 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_47 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_46 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X515 VSS iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=1.27 ps=4.54 w=1 l=0.15
X516 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X517 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_40 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_39 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X518 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X519 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X520 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X521 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X522 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_30 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_29 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X523 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_22 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_21 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X524 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_56 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_57 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X525 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X526 C2_3x7_2.bottom C2_3x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X527 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X528 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 C3_1x5_3.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X529 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_34 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_35 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X530 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_70 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_69 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X531 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_20 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_21 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X532 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_56 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_55 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X533 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X534 VDD iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X535 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X536 C3_1x5_3.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X537 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X538 C3_1x5_3.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl C3_1x5_3.bottom VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X539 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_136 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X540 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_122 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_123 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X541 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_91 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_90 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X542 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_129 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_130 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X543 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_122 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_123 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X544 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X545 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X546 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_81 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_80 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X547 C2_3x7_2.top C2_3x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X548 iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X549 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X550 C3_1x5_3.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X551 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_74 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_73 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X552 C3_1x5_3.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n C3_1x5_3.bottom VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X553 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_37 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_38 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X554 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_113 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_112 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X555 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X556 VSS iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X557 iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X558 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout C3_1x5_3.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X559 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_106 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_105 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X560 iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X561 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X562 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_27 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_28 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X563 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X564 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_83 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_84 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X565 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X566 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_20 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_21 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X567 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X568 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_24 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_25 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X569 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X570 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X571 VSS VDD iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X572 C3_1x5_1.top C3_1x5_1.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X573 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X574 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X575 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_52 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_53 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X576 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_52 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_51 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X577 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_86 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_87 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X578 VDD iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=3.81 ps=8.54 w=3 l=0.15
X579 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_38 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_37 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X580 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_72 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_73 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X581 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X582 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_126 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_127 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X583 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X584 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X585 VDD di_LO_QX iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X586 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X587 VSS iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X588 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X589 VDD iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X590 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X591 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X592 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 C3_1x5_1.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X593 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n di_afe_en VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X594 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X595 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X596 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_121 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_120 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X597 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X598 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X599 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_61 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_62 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X600 VDD iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X601 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_54 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_55 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X602 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X603 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X604 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X605 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X606 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_86 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_87 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X607 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_103 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_104 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X608 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_136 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_135 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X609 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X610 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_2 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_1 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X611 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_19 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_18 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X612 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_76 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_77 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X613 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X614 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_101 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_100 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X615 C2_3x7_2.bottom C2_3x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X616 C3_1x5_3.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X617 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X618 C2_3x7_2.bottom C2_3x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X619 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 C3_1x5_1.top C3_1x5_1.bottom VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X620 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X621 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_113 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_114 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X622 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_51 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_50 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X623 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X624 C2_3x7_2.top C2_3x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X625 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_44 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_43 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X626 C3_1x5_1.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl C3_1x5_1.bottom VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X627 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X628 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X629 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X630 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X631 C3_1x5_3.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X632 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X633 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_34 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_33 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X634 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X635 C3_1x5_3.bottom C3_1x5_3.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X636 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X637 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X638 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X639 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X640 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X641 C2_3x7_2.top C2_3x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X642 C3_1x5_1.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n C3_1x5_1.bottom VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X643 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X644 di_LO_QX VSS iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0.495 ps=3.33 w=3 l=0.15
X645 VDD iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X646 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X647 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X648 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X649 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_59 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_60 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X650 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_85 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_84 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X651 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X652 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X653 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0 ps=0 w=3 l=1
X654 VSS iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X655 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X656 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_116 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_117 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X657 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_133 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_134 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X658 VDD di_afe_en iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X659 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_23 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_24 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X660 C3_1x5_3.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X661 VDD iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=3.81 ps=8.54 w=3 l=0.15
X662 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_59 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_58 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X663 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_75 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_74 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X664 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X665 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X666 VSS iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X667 VDD iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X668 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_68 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_67 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X669 VDD iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X670 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X671 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X672 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_103 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_104 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X673 VDD iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X674 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_31 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_32 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X675 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X676 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_107 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_106 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X677 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_125 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_126 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X678 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin di_LO_QX VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X679 VDD iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X680 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X681 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_84 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_83 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X682 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_100 C2_3x7_2.top VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X683 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X684 C3_1x5_3.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X685 VDD iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X686 iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X687 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_21 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_22 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X688 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_14 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_15 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X689 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X690 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X691 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X692 VSS iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X693 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X694 VSS di_LO_Q iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X695 C3_1x5_1.bottom C3_1x5_1.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X696 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_46 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_47 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X697 VSS VDD iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X698 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X699 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X700 VDD iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X701 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X702 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X703 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X704 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_77 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_76 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X705 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_41 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_42 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X706 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_63 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_62 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X707 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_27 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_28 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X708 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X709 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin di_LO_Q VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X710 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_115 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_114 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X711 vinn_I iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_0 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X712 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X713 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X714 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 C3_1x5_3.top C3_1x5_3.bottom VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X715 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X716 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_89 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_90 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X717 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_41 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_40 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X718 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X719 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_75 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_76 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X720 di_LO_QX VDD iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X721 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n C3_1x5_3.bottom VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X722 VSS VDD iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X723 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_129 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_130 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X724 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_115 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_116 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X725 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X726 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X727 VDD iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X728 C2_3x7_2.top C2_3x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X729 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_97 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_98 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X730 VSS VDD iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X731 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_129 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_128 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X732 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X733 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X734 iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X735 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X736 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_100 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_101 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X737 C3_1x5_3.top C3_1x5_3.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X738 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_90 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_91 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X739 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X740 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_130 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_129 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X741 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X742 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X743 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_13 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_12 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X744 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X745 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X746 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl C3_1x5_3.bottom VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X747 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 C3_1x5_1.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X748 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X749 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X750 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_114 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_113 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X751 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_80 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_81 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X752 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X753 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_45 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_44 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X754 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X755 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X756 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X757 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X758 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout C3_1x5_1.bottom VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X759 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_38 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_37 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X760 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_112 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_113 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X761 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X762 VDD iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X763 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X764 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X765 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X766 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X767 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X768 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X769 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X770 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X771 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_28 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_27 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X772 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X773 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n C3_1x5_1.bottom VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X774 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X775 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X776 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X777 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X778 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_79 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_80 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X779 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_45 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_44 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X780 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_31 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_30 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X781 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout C3_1x5_1.bottom VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X782 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X783 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_60 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_59 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X784 C2_3x7_2.bottom C2_3x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X785 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_93 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_92 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X786 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_43 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_44 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X787 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_79 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_78 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X788 iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X789 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_133 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_132 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X790 VDD iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X791 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_24 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_23 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X792 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_58 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_59 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X793 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl C3_1x5_1.bottom VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X794 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X795 VDD iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X796 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_127 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_128 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X797 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X798 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X799 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_104 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_103 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X800 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X801 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_120 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_121 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X802 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X803 VSS di_afe_en iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X804 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X805 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_126 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_125 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X806 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_62 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_61 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X807 VDD iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X808 VDD iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X809 C2_3x7_2.top C2_3x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X810 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X811 VDD iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X812 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout C3_1x5_3.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X813 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X814 iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X815 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X816 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X817 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X818 C3_1x5_3.bottom C3_1x5_3.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X819 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_104 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_103 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X820 iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X821 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X822 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_63 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_64 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X823 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n C3_1x5_3.bottom VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X824 C1_5x7_2.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_16 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X825 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_3 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_2 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X826 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VDD di_LO_I VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X827 iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X828 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_18 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_19 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X829 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X830 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X831 C3_1x5_1.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X832 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_97 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_96 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X833 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_95 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_96 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X834 C3_1x5_1.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl C3_1x5_1.bottom VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X835 VSS iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X836 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X837 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_50 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_51 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X838 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X839 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_42 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_41 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X840 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X841 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X842 VDD iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=3.81 ps=8.54 w=3 l=0.15
X843 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X844 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_28 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_27 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X845 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_76 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_77 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X846 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_11 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_10 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X847 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_62 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_63 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X848 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl C3_1x5_3.bottom VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X849 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 C3_1x5_1.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X850 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X851 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X852 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X853 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_90 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_89 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X854 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_40 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_41 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X855 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_76 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_75 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X856 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X857 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X858 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X859 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_130 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_129 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X860 C3_1x5_1.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X861 C2_3x7_2.bottom C2_3x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X862 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_116 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_115 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X863 C3_1x5_1.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n C3_1x5_1.bottom VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X864 C3_1x5_1.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X865 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X866 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X867 VSS iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X868 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X869 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X870 C3_1x5_1.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X871 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X872 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_128 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_129 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X873 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X874 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 C3_1x5_3.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X875 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_91 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_92 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X876 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X877 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X878 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n C3_1x5_3.bottom VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X879 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X880 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_84 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_85 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X881 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X882 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_7 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_6 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X883 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_7 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_6 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X884 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X885 iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X886 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X887 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X888 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X889 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_134 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_133 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X890 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X891 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout C3_1x5_3.bottom VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X892 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X893 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_74 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_75 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X894 C2_3x7_2.top C2_3x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X895 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_55 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_54 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X896 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_19 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_20 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X897 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X898 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl C3_1x5_3.bottom VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X899 VSS iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X900 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_32 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_31 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X901 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X902 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_106 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_107 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X903 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_125 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_126 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X904 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X905 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_44 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_45 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X906 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X907 VDD iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X908 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_30 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_31 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X909 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_80 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_79 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X910 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X911 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_22 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_21 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X912 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X913 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X914 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X915 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X916 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X917 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_92 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_93 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X918 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_44 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_43 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X919 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_78 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_79 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X920 C3_1x5_1.top C3_1x5_1.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X921 VSS di_LO_QX iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X922 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X923 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_132 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_133 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X924 vinn_Q iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_0 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X925 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X926 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X927 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X928 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_23 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_24 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X929 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X930 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_121 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_122 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X931 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X932 C3_1x5_1.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X933 C3_1x5_3.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X934 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_114 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_115 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X935 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_0 vinp_Q VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X936 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout C3_1x5_1.bottom VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X937 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X938 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X939 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X940 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_37 C2_3x7_2.bottom VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X941 VSS iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X942 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X943 VDD iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X944 VSS iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X945 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X946 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X947 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_16 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X948 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_98 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_97 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X949 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_2 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_3 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X950 C3_1x5_1.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X951 C3_1x5_3.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X952 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X953 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_57 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_58 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X954 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X955 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X956 VSS VDD iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X957 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X958 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X959 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_96 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_97 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X960 iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X961 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_12 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_13 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X962 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_89 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_90 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X963 di_LO_Q VSS iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0.495 ps=3.33 w=3 l=0.15
X964 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X965 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X966 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X967 C2_3x7_2.bottom C2_3x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X968 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X969 VDD iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X970 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X971 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_44 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_45 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X972 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_5 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_4 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X973 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X974 VSS iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X975 C2_3x7_2.top C2_3x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X976 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X977 C3_1x5_1.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X978 C3_1x5_3.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X979 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X980 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X981 VSS iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=1.27 ps=4.54 w=1 l=0.15
X982 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X983 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X984 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X985 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X986 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X987 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X988 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X989 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X990 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X991 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X992 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X993 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X994 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_65 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_66 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X995 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X996 C2_3x7_2.top C2_3x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X997 C3_1x5_1.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X998 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X999 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 C3_1x5_1.top C3_1x5_1.bottom VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1000 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_6 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_7 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1001 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1002 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_119 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_118 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1003 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1004 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 C3_1x5_3.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1005 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_20 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_19 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1006 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1007 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_128 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_127 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1008 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_54 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_55 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1009 VSS iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1010 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1011 VDD iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1012 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1013 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1014 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1015 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_119 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_120 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1016 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 C3_1x5_1.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1017 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1018 C3_1x5_3.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1019 VSS iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1020 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1021 VSS iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1022 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_71 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_70 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1023 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1024 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n C3_1x5_1.bottom VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1025 di_LO_Q VDD iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X1026 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_64 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_63 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1027 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_0 vinp_I VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1028 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1029 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1030 VSS iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1031 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1032 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1033 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1034 VDD di_afe_en iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1035 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1036 VDD iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X1037 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_96 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_95 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1038 C3_1x5_3.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1039 VDD iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1040 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_18 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1041 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_83 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_82 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1042 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_47 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_48 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1043 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1044 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_69 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_68 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1045 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_33 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_34 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1046 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1047 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1048 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1049 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_10 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_11 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1050 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl C3_1x5_1.bottom VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1051 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1052 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout C3_1x5_3.bottom VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1053 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin di_LO_I VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1054 di_LO_I VSS iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0.495 ps=3.33 w=3 l=0.15
X1055 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1056 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1057 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_95 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_96 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1058 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_135 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_136 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1059 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1060 VSS iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1061 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1062 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1063 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_37 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1064 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1065 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1066 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1067 C3_1x5_1.bottom C3_1x5_1.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1068 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1069 C2_3x7_2.top C2_3x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1070 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_92 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_91 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1071 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1072 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1073 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1074 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=0 ps=0 w=9 l=1
X1075 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1076 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 C3_1x5_1.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1077 iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1078 C3_1x5_3.top C3_1x5_3.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1079 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1080 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout C3_1x5_3.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1081 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_6 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_7 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1082 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1083 iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1084 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1085 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_93 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_94 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1086 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1087 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1088 VSS VDD iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X1089 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_5 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_6 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1090 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1091 VDD iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1092 iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1093 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_126 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_125 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1094 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1095 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_9 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_8 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1096 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1097 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1098 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1099 C2_3x7_2.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_100 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1100 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_83 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_84 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1101 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_85 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_86 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1102 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_51 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_50 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1103 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1104 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1105 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1106 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1107 VDD iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1108 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1109 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1110 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_41 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_40 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1111 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_66 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_65 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1112 C3_1x5_1.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_98 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1113 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1114 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X1115 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1116 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout C3_1x5_1.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1117 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 C3_1x5_3.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1118 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1119 C2_3x7_2.bottom C2_3x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1120 iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1121 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_118 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_119 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1122 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1123 VSS VDD iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X1124 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n C3_1x5_1.bottom VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1125 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_24 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_23 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1126 iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1127 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VDD di_LO_IX VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X1128 C3_1x5_1.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1129 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1130 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_122 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_121 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1131 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1132 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1133 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1134 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 C3_1x5_3.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1135 iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1136 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_9 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_10 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1137 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1138 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl C3_1x5_1.bottom VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1139 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout C3_1x5_3.bottom VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1140 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1141 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout C3_1x5_1.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1142 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_123 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_124 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1143 VDD di_afe_en iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1144 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_57 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_58 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1145 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_23 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_22 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1146 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_9 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_8 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1147 VDD iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1148 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_65 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_64 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1149 VDD iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1150 VDD iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1151 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout C3_1x5_1.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1152 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1153 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_58 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_57 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1154 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_103 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_102 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1155 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1156 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1157 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1158 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1159 C2_3x7_2.bottom C2_3x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1160 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_48 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_47 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1161 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_34 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_33 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1162 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_82 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_83 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1163 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_90 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_89 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1164 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1165 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1166 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_68 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_69 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1167 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n C3_1x5_1.bottom VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1168 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_11 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_12 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1169 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1170 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1171 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1172 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 C3_1x5_3.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1173 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_96 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_95 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1174 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_4 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_5 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1175 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_136 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_135 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1176 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1177 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1178 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin di_LO_I VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1179 C3_1x5_1.bottom C3_1x5_1.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1180 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1181 C2_3x7_2.bottom C2_3x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1182 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_53 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_54 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1183 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1184 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl C3_1x5_1.bottom VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1185 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1186 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1187 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1188 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1189 VSS di_afe_en iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1190 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1191 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_27 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_26 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1192 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_61 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_62 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1193 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_13 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_12 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1194 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n C3_1x5_3.bottom VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1195 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1196 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1197 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 C3_1x5_3.top C3_1x5_3.bottom VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1198 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1199 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_39 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_40 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1200 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_61 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_60 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1201 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_25 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_26 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1202 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_55 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_56 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1203 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_136 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1204 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout C3_1x5_3.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1205 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_115 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_114 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1206 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1207 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout C3_1x5_3.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1208 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_6 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_5 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1209 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1210 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1211 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1212 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_87 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_88 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1213 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1214 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl C3_1x5_3.bottom VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1215 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_50 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_51 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1216 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_100 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1217 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1218 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_86 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_85 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1219 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_120 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_119 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1220 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_3 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_2 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1221 VSS iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=1.27 ps=4.54 w=1 l=0.15
X1222 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_77 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_78 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1223 C3_1x5_1.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1224 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1225 VSS iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1226 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_98 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1227 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_70 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_71 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1228 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n di_afe_en VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1229 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1230 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1231 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_35 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_34 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1232 VSS iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1233 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n di_afe_en VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1234 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1235 VSS iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1236 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1237 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1238 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1239 VDD di_LO_Q iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1240 C3_1x5_1.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1241 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1242 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1243 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1244 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_18 C1_5x7_2.top VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1245 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1246 C2_3x7_2.top C2_3x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1247 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1248 iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1249 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin di_LO_Q VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1250 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1251 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1252 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_10 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_9 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1253 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_43 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_42 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1254 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1255 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1256 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1257 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1258 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1259 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1260 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_22 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_23 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1261 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_8 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_9 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1262 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_58 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_57 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1263 VDD iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=3.81 ps=8.54 w=3 l=0.15
X1264 VDD di_LO_I iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1265 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_79 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_78 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1266 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_117 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_118 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1267 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1268 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 C3_1x5_1.top C3_1x5_1.bottom VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1269 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1270 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_102 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_103 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1271 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1272 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_111 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_110 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1273 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_69 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_68 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1274 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1275 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_25 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_26 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1276 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_101 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_100 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1277 C2_3x7_2.bottom C2_3x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1278 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1279 VDD iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1280 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1281 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1282 C3_1x5_3.bottom C3_1x5_3.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1283 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_94 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_93 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1284 VSS iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1285 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1286 C3_1x5_3.bottom C3_1x5_3.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1287 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_15 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_16 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1288 C2_3x7_2.top C2_3x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1289 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_2 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1290 VDD iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X1291 iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1292 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1293 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1294 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_8 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_9 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1295 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1296 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1297 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1298 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_84 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_83 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1299 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1300 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1301 VSS iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1302 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1303 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_47 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_48 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1304 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1305 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1306 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_40 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_41 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1307 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1308 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X1309 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_26 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_27 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1310 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_62 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_61 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1311 VSS di_afe_en iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1312 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1313 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1314 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_12 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_13 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1315 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1316 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1317 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1318 C3_1x5_1.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1319 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1320 VSS iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1321 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1322 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_40 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_39 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1323 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1324 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_26 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_25 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1325 C2_3x7_2.bottom C2_3x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1326 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_60 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_61 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1327 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n di_afe_en VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1328 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_114 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_115 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1329 VDD iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1330 VSS iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1331 VSS iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1332 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1333 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1334 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1335 C3_1x5_1.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1336 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1337 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_81 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_82 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1338 VDD iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1339 iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1340 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_131 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_130 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1341 di_LO_IX VSS iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0.495 ps=3.33 w=3 l=0.15
X1342 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_71 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_72 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1343 iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1344 C3_1x5_1.bottom C3_1x5_1.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1345 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_124 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_123 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1346 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1347 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1348 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_64 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_65 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1349 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_49 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_48 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1350 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1351 VDD iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1352 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1353 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1354 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1355 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_39 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_38 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1356 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1357 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_89 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_88 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1358 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_53 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_54 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1359 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1360 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 C3_1x5_3.top C3_1x5_3.bottom VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1361 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_12 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_11 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1362 iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1363 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1364 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1365 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n C3_1x5_3.bottom VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1366 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1367 VDD iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X1368 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_42 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_43 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1369 VSS VDD iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X1370 VDD iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1371 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1372 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1373 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1374 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_54 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_53 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1375 iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1376 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1377 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1378 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1379 C3_1x5_3.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1380 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1381 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_73 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_72 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1382 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 C3_1x5_1.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1383 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X1384 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl C3_1x5_3.bottom VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1385 C2_3x7_2.top C2_3x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1386 VSS di_LO_I iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1387 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1388 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1389 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_105 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_104 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1390 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_63 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_62 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1391 C3_1x5_3.top C3_1x5_3.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1392 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout C3_1x5_1.bottom VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1393 VSS VDD iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X1394 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1395 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1396 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_56 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_55 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1397 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1398 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1399 VSS VDD iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X1400 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_136 C3_1x5_3.bottom VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1401 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_107 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_106 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1402 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1403 C3_1x5_3.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1404 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_19 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_20 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1405 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_95 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_94 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1406 VSS VDD iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X1407 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout C3_1x5_1.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1408 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1409 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1410 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1411 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1412 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_88 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_87 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1413 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_2 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_1 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1414 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1415 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_105 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_106 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1416 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_9 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_10 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1417 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_51 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_52 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1418 VDD di_afe_en iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1419 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout C3_1x5_1.bottom VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1420 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1421 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1422 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_2 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_3 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1423 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1424 C3_1x5_3.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1425 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_78 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_77 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1426 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_41 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_42 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1427 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1428 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1429 VSS iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1430 VSS VDD iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X1431 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_34 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_35 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1432 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1433 C3_1x5_1.top C3_1x5_1.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1434 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1435 C2_3x7_2.bottom C2_3x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1436 VDD iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1437 VDD iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1438 VDD iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1439 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1440 C3_1x5_3.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1441 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1442 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1443 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1444 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1445 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1446 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_29 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_30 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1447 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_65 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_64 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1448 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_15 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_16 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1449 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_135 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_134 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1450 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n di_afe_en VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1451 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1452 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1453 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1454 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1455 VSS VDD iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X1456 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_109 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_110 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1457 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_29 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_28 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1458 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_85 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_86 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1459 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_63 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_64 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1460 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_125 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_124 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1461 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_131 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_132 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1462 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n C3_1x5_3.bottom VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1463 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1464 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_117 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_118 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1465 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_78 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_79 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1466 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_118 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_117 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1467 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_43 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_42 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1468 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_0 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1469 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_109 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_108 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1470 iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1471 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_68 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_69 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1472 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_54 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_53 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1473 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_110 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_111 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1474 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_88 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_89 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1475 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 C3_1x5_1.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1476 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_33 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_32 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1477 C2_3x7_2.bottom C2_3x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1478 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl C3_1x5_3.bottom VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1479 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 C3_1x5_1.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1480 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_26 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_25 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1481 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_100 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_101 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1482 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n C3_1x5_1.bottom VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1483 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1484 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1485 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1486 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1487 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1488 VSS iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1489 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1490 iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1491 C3_1x5_1.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1492 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_16 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_15 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1493 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1494 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1495 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1496 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1497 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1498 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1499 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1500 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_48 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_47 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1501 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1502 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl C3_1x5_1.bottom VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1503 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1504 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_47 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_46 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1505 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_81 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_82 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1506 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_33 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_32 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1507 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1508 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_67 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_68 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1509 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_19 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_18 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1510 C2_3x7_2.top C2_3x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1511 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1512 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_121 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_122 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1513 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_67 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_66 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1514 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1515 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1516 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout C3_1x5_3.bottom VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1517 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1518 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1519 iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1520 VSS iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1521 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_45 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_46 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1522 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X1523 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1524 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_115 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_116 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1525 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1526 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_135 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_134 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1527 C3_1x5_3.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1528 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_57 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_56 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1529 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_121 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_120 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1530 C3_1x5_3.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl C3_1x5_3.bottom VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1531 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_106 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_107 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1532 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_109 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_108 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1533 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1534 VSS iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1535 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1536 VSS VDD iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X1537 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_106 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_105 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1538 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_82 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_81 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1539 C3_1x5_3.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl C3_1x5_3.bottom VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1540 C3_1x5_3.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1541 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1542 C3_1x5_3.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n C3_1x5_3.bottom VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1543 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_130 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_131 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1544 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_72 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_71 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1545 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1546 iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1547 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_48 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_49 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1548 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1549 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1550 C3_1x5_3.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n C3_1x5_3.bottom VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1551 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_5 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_4 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1552 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1553 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout C3_1x5_1.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1554 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_38 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_39 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1555 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 C3_1x5_1.top C3_1x5_1.bottom VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1556 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1557 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_49 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_50 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1558 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_85 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_84 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1559 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1560 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1561 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 C3_1x5_3.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1562 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1563 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1564 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1565 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1566 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_30 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_29 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1567 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_64 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_65 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1568 C2_3x7_2.top C2_3x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1569 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_16 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_15 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1570 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_49 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_48 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1571 VSS iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1572 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1573 VSS iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1574 iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1575 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X1576 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout C3_1x5_1.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1577 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_110 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_109 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1578 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n C3_1x5_3.bottom VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1579 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_28 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_29 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1580 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_64 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_63 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1581 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_132 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_131 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1582 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_118 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_117 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1583 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1584 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1585 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_79 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_80 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1586 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1587 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1588 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_108 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_109 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1589 iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1590 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1591 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_72 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_73 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1592 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1593 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_37 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1594 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1595 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_111 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_112 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1596 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1597 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1598 VSS VDD iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X1599 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1600 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl C3_1x5_3.bottom VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1601 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_104 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_105 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1602 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_62 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_63 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1603 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_27 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_26 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1604 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1605 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1606 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1607 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_20 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_19 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1608 VSS di_LO_IX iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1609 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_94 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_95 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1610 C2_3x7_2.bottom C2_3x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1611 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_7 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_8 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1612 C3_1x5_3.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1613 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1614 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_52 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_51 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1615 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_10 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_9 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1616 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin di_LO_IX VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1617 iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1618 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1619 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1620 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1621 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1622 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1623 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_46 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_47 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1624 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_82 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_81 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1625 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1626 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_32 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_33 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1627 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_68 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_67 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1628 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_42 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_41 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1629 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1630 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_18 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_19 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1631 VDD iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X1632 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_122 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_121 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1633 C3_1x5_3.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1634 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1635 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1636 iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1637 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1638 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 C3_1x5_3.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1639 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1640 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1641 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_46 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_45 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1642 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1643 VDD iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X1644 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1645 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_134 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_135 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1646 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_120 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_121 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1647 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1648 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X1649 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1650 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1651 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1652 C2_3x7_2.bottom C2_3x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1653 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1654 VDD iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1655 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1656 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 C3_1x5_1.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1657 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_103 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_102 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1658 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1659 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1660 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1661 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X1662 VDD iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1663 C3_1x5_3.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1664 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_134 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_135 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1665 iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1666 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1667 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1668 VDD iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1669 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_86 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_85 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1670 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n C3_1x5_1.bottom VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1671 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_124 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_125 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1672 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1673 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_49 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_50 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1674 VSS VDD iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X1675 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1676 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1677 iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1678 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout C3_1x5_3.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1679 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_42 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_43 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1680 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_0 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_1 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1681 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 C3_1x5_3.top C3_1x5_3.bottom VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1682 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_4 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_5 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1683 iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1684 C3_1x5_3.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1685 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.93 pd=6.62 as=0 ps=0 w=3 l=0.15
X1686 C3_1x5_1.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n vout_RF VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1687 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1688 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_50 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_49 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1689 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_84 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_85 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1690 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_32 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_33 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1691 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VDD VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1692 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl C3_1x5_1.bottom VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1693 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1694 VDD iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X1695 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1696 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout C3_1x5_3.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1697 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1698 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_48 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_49 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1699 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1700 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1701 VDD iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1702 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1703 C1_5x7_2.top C1_5x7_2.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1704 C3_1x5_1.bottom iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1705 C2_3x7_2.bottom C2_3x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1706 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1707 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 C3_1x5_1.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1708 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1709 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_133 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_132 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1710 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout C3_1x5_3.top iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1711 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1712 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1713 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n C3_1x5_3.bottom VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1714 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_66 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_67 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1715 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl vout_RF VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1716 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1717 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0 ps=0 w=3 l=1
X1718 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1719 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_116 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_115 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1720 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1721 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_113 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_112 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1722 VDD iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1723 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_56 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_57 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1724 C3_1x5_3.top C3_1x5_3.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1725 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1726 iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1727 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1728 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_108 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_109 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1729 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_8 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_7 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1730 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_31 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_30 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1731 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl C3_1x5_3.bottom VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1732 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1733 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1734 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1735 C1_5x7_2.bottom C1_5x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1736 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_59 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_58 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1737 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 C3_1x5_3.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1738 VDD iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=3.81 ps=8.54 w=3 l=0.15
X1739 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1740 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1741 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0 ps=0 w=3 l=0.15
X1742 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1743 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1744 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1745 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1746 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n di_afe_en VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1747 C3_1x5_1.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1748 vout_RF iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n C3_1x5_1.bottom VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1749 C3_1x5_1.top C3_1x5_1.bottom sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1750 vout_RF iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1751 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1752 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_5 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_6 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1753 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_71 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_72 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1754 C2_3x7_2.bottom C2_3x7_2.top sky130_fd_pr__cap_mim_m3_1 l=3 w=3
X1755 VDD iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VDD sky130_fd_pr__pfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1756 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 C3_1x5_3.bottom iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1757 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VDD sky130_fd_pr__pfet_01v8_lvt ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1758 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_35 C2_3x7_2.bottom VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1759 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0 ps=0 w=1 l=0.15
X1760 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_71 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_70 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1761 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_125 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_124 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1762 VSS iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=1.27 ps=4.54 w=1 l=0.15
X1763 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_97 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_96 VSS sky130_fd_pr__res_xhigh_po_0p35 l=2
C0 vinn_Q VSS 3.84856f
C1 di_LO_Q VSS 4.18304f
C2 di_LO_QX VSS 4.18304f
C3 vinp_Q VSS 3.84856f
C4 vinn_I VSS 3.84856f
C5 di_LO_I VSS 4.18304f
C6 vout_RF VSS 64.6665f
C7 di_afe_en VSS 16.084f
C8 di_LO_IX VSS 4.18304f
C9 vinp_I VSS 3.84856f
C10 VDD VSS 1.18296p
C11 iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VSS 11.5065f
C12 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VSS 4.48926f
C13 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VSS 2.83622f
C14 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_136 VSS 1.22562f
C15 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_135 VSS 1.22562f
C16 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_134 VSS 1.22562f
C17 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_133 VSS 1.22629f
C18 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_132 VSS 1.22562f
C19 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_131 VSS 1.22762f
C20 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_130 VSS 1.22562f
C21 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_129 VSS 1.22562f
C22 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_128 VSS 1.22629f
C23 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_127 VSS 1.22696f
C24 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_126 VSS 1.22562f
C25 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_125 VSS 1.22562f
C26 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_124 VSS 1.22562f
C27 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_123 VSS 1.22629f
C28 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_122 VSS 1.22696f
C29 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_121 VSS 1.22762f
C30 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_120 VSS 1.22562f
C31 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_119 VSS 1.22562f
C32 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_118 VSS 1.22562f
C33 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_117 VSS 1.22696f
C34 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_116 VSS 1.22562f
C35 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_115 VSS 1.22562f
C36 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_114 VSS 1.22562f
C37 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_113 VSS 1.22629f
C38 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_112 VSS 1.22562f
C39 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_111 VSS 1.22762f
C40 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_110 VSS 1.22562f
C41 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_109 VSS 1.22562f
C42 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_108 VSS 1.22629f
C43 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_107 VSS 1.22696f
C44 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_106 VSS 1.22762f
C45 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_105 VSS 1.22562f
C46 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_104 VSS 1.22562f
C47 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_103 VSS 1.22629f
C48 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_102 VSS 1.22696f
C49 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_101 VSS 1.22762f
C50 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_100 VSS 1.22562f
C51 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_98 VSS 1.22629f
C52 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_97 VSS 1.22696f
C53 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_96 VSS 1.22562f
C54 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_95 VSS 1.22562f
C55 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_94 VSS 1.22562f
C56 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_93 VSS 1.22629f
C57 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_92 VSS 1.22696f
C58 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_91 VSS 1.22762f
C59 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_90 VSS 1.22562f
C60 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_89 VSS 1.22562f
C61 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_88 VSS 1.22562f
C62 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_87 VSS 1.22696f
C63 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_86 VSS 1.22562f
C64 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_85 VSS 1.22562f
C65 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_84 VSS 1.22562f
C66 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_83 VSS 1.22629f
C67 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_82 VSS 1.22696f
C68 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_81 VSS 1.22762f
C69 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_80 VSS 1.22562f
C70 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_79 VSS 1.22562f
C71 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_78 VSS 1.22629f
C72 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_77 VSS 1.22696f
C73 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_76 VSS 1.22562f
C74 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_75 VSS 1.22562f
C75 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_74 VSS 1.22562f
C76 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_73 VSS 1.22629f
C77 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_72 VSS 1.22696f
C78 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_71 VSS 1.22562f
C79 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_70 VSS 1.22562f
C80 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_69 VSS 1.22562f
C81 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_68 VSS 1.22629f
C82 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_67 VSS 1.22696f
C83 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_66 VSS 1.22762f
C84 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_65 VSS 1.22562f
C85 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_64 VSS 1.22562f
C86 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_63 VSS 1.22629f
C87 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_62 VSS 1.22696f
C88 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_61 VSS 1.22762f
C89 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_60 VSS 1.22562f
C90 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_59 VSS 1.22562f
C91 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_58 VSS 1.22629f
C92 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_57 VSS 1.22562f
C93 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_56 VSS 1.22762f
C94 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_55 VSS 1.22562f
C95 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_54 VSS 1.22562f
C96 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_53 VSS 1.22629f
C97 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_52 VSS 1.22696f
C98 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_51 VSS 1.22762f
C99 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_50 VSS 1.22562f
C100 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_49 VSS 1.22562f
C101 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_48 VSS 1.22629f
C102 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_47 VSS 1.22696f
C103 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_46 VSS 1.22562f
C104 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_45 VSS 1.22562f
C105 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_44 VSS 1.22562f
C106 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_43 VSS 1.22629f
C107 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_42 VSS 1.22696f
C108 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_41 VSS 1.22762f
C109 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_40 VSS 1.22562f
C110 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_39 VSS 1.22562f
C111 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_38 VSS 1.22629f
C112 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_37 VSS 1.22696f
C113 C2_3x7_2.bottom VSS 56.048f
C114 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_35 VSS 1.22829f
C115 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_34 VSS 1.22562f
C116 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_33 VSS 1.22629f
C117 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_32 VSS 1.22696f
C118 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_31 VSS 1.22762f
C119 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_30 VSS 1.22562f
C120 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_29 VSS 1.22562f
C121 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_28 VSS 1.22629f
C122 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_27 VSS 1.22696f
C123 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_26 VSS 1.22562f
C124 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_25 VSS 1.22562f
C125 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_24 VSS 1.22562f
C126 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_23 VSS 1.22629f
C127 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_22 VSS 1.22696f
C128 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_21 VSS 1.22762f
C129 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_20 VSS 1.22562f
C130 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_19 VSS 1.22562f
C131 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_18 VSS 1.22629f
C132 C1_5x7_2.bottom VSS 78.81621f
C133 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_16 VSS 1.22562f
C134 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_15 VSS 1.22562f
C135 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_14 VSS 1.22562f
C136 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_13 VSS 1.22629f
C137 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_12 VSS 1.22562f
C138 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_11 VSS 1.22762f
C139 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_10 VSS 1.22562f
C140 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_9 VSS 1.22562f
C141 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_8 VSS 1.22629f
C142 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_7 VSS 1.22696f
C143 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_6 VSS 1.22562f
C144 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_5 VSS 1.22562f
C145 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_4 VSS 1.22562f
C146 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_3 VSS 1.22629f
C147 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_2 VSS 1.22896f
C148 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_1 VSS 1.22562f
C149 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_0 VSS 1.22562f
C150 iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VSS 14.3155f
C151 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VSS 4.48926f
C152 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VSS 7.66312f
C153 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VSS 7.89561f
C154 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin VSS 2.82434f
C155 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS 3.36642f
C156 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS 3.36642f
C157 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VSS 2.49069f
C158 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS 3.36642f
C159 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS 3.36642f
C160 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS 3.36642f
C161 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS 3.36642f
C162 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS 3.36642f
C163 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VSS 2.49069f
C164 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS 3.36642f
C165 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS 3.36642f
C166 iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VSS 11.5086f
C167 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VSS 4.48926f
C168 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VSS 2.83622f
C169 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VSS 7.84314f
C170 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VSS 7.84314f
C171 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VSS 5.82216f
C172 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VSS 7.84314f
C173 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VSS 51.5669f
C174 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VSS 7.84314f
C175 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VSS 7.84314f
C176 C3_1x5_1.bottom VSS 71.3916f
C177 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VSS 7.84314f
C178 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VSS 7.84314f
C179 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VSS 5.82216f
C180 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VSS 7.84314f
C181 C3_1x5_1.top VSS 33.3927f
C182 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS 75.0436f
C183 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VSS 7.84314f
C184 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VSS 37.237f
C185 iq_modulator_half_1.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VSS 14.3155f
C186 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VSS 4.48926f
C187 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VSS 7.66312f
C188 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VSS 7.89561f
C189 iq_modulator_half_1.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin VSS 2.82434f
C190 C3_1x5_3.bottom VSS 77.9315f
C191 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_136 VSS 1.22562f
C192 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_135 VSS 1.22562f
C193 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_134 VSS 1.22562f
C194 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_133 VSS 1.22562f
C195 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_132 VSS 1.22696f
C196 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_131 VSS 1.22562f
C197 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_130 VSS 1.22562f
C198 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_129 VSS 1.22562f
C199 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_128 VSS 1.22629f
C200 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_127 VSS 1.22562f
C201 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_126 VSS 1.22562f
C202 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_125 VSS 1.22562f
C203 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_124 VSS 1.22562f
C204 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_123 VSS 1.22629f
C205 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_122 VSS 1.22696f
C206 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_121 VSS 1.22562f
C207 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_120 VSS 1.22562f
C208 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_119 VSS 1.22629f
C209 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_118 VSS 1.22629f
C210 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_117 VSS 1.22562f
C211 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_116 VSS 1.22562f
C212 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_115 VSS 1.22562f
C213 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_114 VSS 1.22562f
C214 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_113 VSS 1.22562f
C215 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_112 VSS 1.22696f
C216 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_111 VSS 1.22562f
C217 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_110 VSS 1.22562f
C218 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_109 VSS 1.22562f
C219 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_108 VSS 1.22629f
C220 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_107 VSS 1.22696f
C221 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_106 VSS 1.22562f
C222 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_105 VSS 1.22562f
C223 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_104 VSS 1.22562f
C224 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_103 VSS 1.22629f
C225 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_102 VSS 1.22696f
C226 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_101 VSS 1.22562f
C227 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_100 VSS 1.22562f
C228 C3_1x5_3.top VSS 39.0581f
C229 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_98 VSS 1.22629f
C230 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_97 VSS 1.22562f
C231 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_96 VSS 1.22562f
C232 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_95 VSS 1.22562f
C233 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_94 VSS 1.22562f
C234 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_93 VSS 1.22629f
C235 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_92 VSS 1.22696f
C236 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_91 VSS 1.22562f
C237 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_90 VSS 1.22562f
C238 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_89 VSS 1.22629f
C239 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_88 VSS 1.22629f
C240 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_87 VSS 1.22562f
C241 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_86 VSS 1.22562f
C242 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_85 VSS 1.22562f
C243 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_84 VSS 1.22562f
C244 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_83 VSS 1.22629f
C245 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_82 VSS 1.22696f
C246 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_81 VSS 1.22562f
C247 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_80 VSS 1.22562f
C248 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_79 VSS 1.22562f
C249 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_78 VSS 1.22629f
C250 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_77 VSS 1.22562f
C251 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_76 VSS 1.22562f
C252 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_75 VSS 1.22562f
C253 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_74 VSS 1.22562f
C254 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_73 VSS 1.22629f
C255 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_72 VSS 1.22562f
C256 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_71 VSS 1.22562f
C257 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_70 VSS 1.22562f
C258 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_69 VSS 1.22562f
C259 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_68 VSS 1.22629f
C260 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_67 VSS 1.22696f
C261 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_66 VSS 1.22562f
C262 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_65 VSS 1.22562f
C263 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_64 VSS 1.22562f
C264 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_63 VSS 1.22629f
C265 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_62 VSS 1.22696f
C266 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_61 VSS 1.22562f
C267 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_60 VSS 1.22562f
C268 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_59 VSS 1.22562f
C269 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_58 VSS 1.22562f
C270 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_57 VSS 1.22696f
C271 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_56 VSS 1.22562f
C272 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_55 VSS 1.22562f
C273 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_54 VSS 1.22562f
C274 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_53 VSS 1.22629f
C275 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_52 VSS 1.22696f
C276 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_51 VSS 1.22562f
C277 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_50 VSS 1.22562f
C278 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_49 VSS 1.22562f
C279 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_48 VSS 1.22629f
C280 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_47 VSS 1.22562f
C281 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_46 VSS 1.22562f
C282 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_45 VSS 1.22562f
C283 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_44 VSS 1.22562f
C284 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_43 VSS 1.22629f
C285 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_42 VSS 1.22696f
C286 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_41 VSS 1.22562f
C287 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_40 VSS 1.22562f
C288 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_39 VSS 1.22562f
C289 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_38 VSS 1.22629f
C290 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_37 VSS 1.22562f
C291 C2_3x7_2.top VSS 59.6624f
C292 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_35 VSS 1.22562f
C293 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_34 VSS 1.22562f
C294 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_33 VSS 1.22629f
C295 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_32 VSS 1.22696f
C296 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_31 VSS 1.22562f
C297 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_30 VSS 1.22562f
C298 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_29 VSS 1.22562f
C299 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_28 VSS 1.22629f
C300 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_27 VSS 1.22562f
C301 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_26 VSS 1.22562f
C302 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_25 VSS 1.22562f
C303 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_24 VSS 1.22562f
C304 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_23 VSS 1.22629f
C305 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_22 VSS 1.22696f
C306 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_21 VSS 1.22562f
C307 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_20 VSS 1.22562f
C308 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_19 VSS 1.22562f
C309 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_18 VSS 1.22629f
C310 C1_5x7_2.top VSS 80.2351f
C311 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_16 VSS 1.22562f
C312 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_15 VSS 1.22562f
C313 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_14 VSS 1.22562f
C314 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_13 VSS 1.22562f
C315 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_12 VSS 1.22696f
C316 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_11 VSS 1.22562f
C317 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_10 VSS 1.22562f
C318 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_9 VSS 1.22562f
C319 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_8 VSS 1.22629f
C320 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_7 VSS 1.22562f
C321 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_6 VSS 1.22562f
C322 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_5 VSS 1.22562f
C323 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_4 VSS 1.22562f
C324 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_3 VSS 1.22896f
C325 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_2 VSS 1.22562f
C326 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_1 VSS 1.22562f
C327 iq_modulator_half_1.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_0 VSS 1.22562f
C328 iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl_n VSS 11.5065f
C329 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_1.vin VSS 4.48926f
C330 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.transmission_gate_wo_dummy_0.v_b VSS 2.83622f
C331 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_136 VSS 1.22562f
C332 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_135 VSS 1.22562f
C333 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_134 VSS 1.22562f
C334 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_133 VSS 1.22629f
C335 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_132 VSS 1.22562f
C336 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_131 VSS 1.22762f
C337 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_130 VSS 1.22562f
C338 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_129 VSS 1.22562f
C339 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_128 VSS 1.22629f
C340 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_127 VSS 1.22696f
C341 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_126 VSS 1.22562f
C342 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_125 VSS 1.22562f
C343 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_124 VSS 1.22562f
C344 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_123 VSS 1.22629f
C345 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_122 VSS 1.22696f
C346 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_121 VSS 1.22762f
C347 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_120 VSS 1.22562f
C348 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_119 VSS 1.22562f
C349 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_118 VSS 1.22562f
C350 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_117 VSS 1.22696f
C351 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_116 VSS 1.22562f
C352 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_115 VSS 1.22562f
C353 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_114 VSS 1.22562f
C354 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_113 VSS 1.22629f
C355 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_112 VSS 1.22562f
C356 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_111 VSS 1.22762f
C357 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_110 VSS 1.22562f
C358 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_109 VSS 1.22562f
C359 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_108 VSS 1.22629f
C360 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_107 VSS 1.22696f
C361 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_106 VSS 1.22762f
C362 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_105 VSS 1.22562f
C363 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_104 VSS 1.22562f
C364 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_103 VSS 1.22629f
C365 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_102 VSS 1.22696f
C366 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_101 VSS 1.22762f
C367 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_100 VSS 1.22562f
C368 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_98 VSS 1.22629f
C369 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_97 VSS 1.22696f
C370 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_96 VSS 1.22562f
C371 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_95 VSS 1.22562f
C372 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_94 VSS 1.22562f
C373 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_93 VSS 1.22629f
C374 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_92 VSS 1.22696f
C375 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_91 VSS 1.22762f
C376 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_90 VSS 1.22562f
C377 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_89 VSS 1.22562f
C378 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_88 VSS 1.22562f
C379 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_87 VSS 1.22696f
C380 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_86 VSS 1.22562f
C381 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_85 VSS 1.22562f
C382 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_84 VSS 1.22562f
C383 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_83 VSS 1.22629f
C384 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_82 VSS 1.22696f
C385 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_81 VSS 1.22762f
C386 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_80 VSS 1.22562f
C387 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_79 VSS 1.22562f
C388 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_78 VSS 1.22629f
C389 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_77 VSS 1.22696f
C390 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_76 VSS 1.22562f
C391 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_75 VSS 1.22562f
C392 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_74 VSS 1.22562f
C393 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_73 VSS 1.22629f
C394 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_72 VSS 1.22696f
C395 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_71 VSS 1.22562f
C396 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_70 VSS 1.22562f
C397 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_69 VSS 1.22562f
C398 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_68 VSS 1.22629f
C399 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_67 VSS 1.22696f
C400 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_66 VSS 1.22762f
C401 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_65 VSS 1.22562f
C402 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_64 VSS 1.22562f
C403 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_63 VSS 1.22629f
C404 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_62 VSS 1.22696f
C405 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_61 VSS 1.22762f
C406 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_60 VSS 1.22562f
C407 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_59 VSS 1.22562f
C408 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_58 VSS 1.22629f
C409 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_57 VSS 1.22562f
C410 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_56 VSS 1.22762f
C411 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_55 VSS 1.22562f
C412 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_54 VSS 1.22562f
C413 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_53 VSS 1.22629f
C414 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_52 VSS 1.22696f
C415 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_51 VSS 1.22762f
C416 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_50 VSS 1.22562f
C417 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_49 VSS 1.22562f
C418 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_48 VSS 1.22629f
C419 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_47 VSS 1.22696f
C420 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_46 VSS 1.22562f
C421 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_45 VSS 1.22562f
C422 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_44 VSS 1.22562f
C423 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_43 VSS 1.22629f
C424 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_42 VSS 1.22696f
C425 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_41 VSS 1.22762f
C426 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_40 VSS 1.22562f
C427 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_39 VSS 1.22562f
C428 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_38 VSS 1.22629f
C429 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_37 VSS 1.22696f
C430 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2n VSS 59.4865f
C431 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_35 VSS 1.22829f
C432 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_34 VSS 1.22562f
C433 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_33 VSS 1.22629f
C434 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_32 VSS 1.22696f
C435 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_31 VSS 1.22762f
C436 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_30 VSS 1.22562f
C437 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_29 VSS 1.22562f
C438 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_28 VSS 1.22629f
C439 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_27 VSS 1.22696f
C440 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_26 VSS 1.22562f
C441 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_25 VSS 1.22562f
C442 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_24 VSS 1.22562f
C443 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_23 VSS 1.22629f
C444 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_22 VSS 1.22696f
C445 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_21 VSS 1.22762f
C446 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_20 VSS 1.22562f
C447 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_19 VSS 1.22562f
C448 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_18 VSS 1.22629f
C449 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1n VSS 79.4888f
C450 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_16 VSS 1.22562f
C451 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_15 VSS 1.22562f
C452 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_14 VSS 1.22562f
C453 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_13 VSS 1.22629f
C454 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_12 VSS 1.22562f
C455 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_11 VSS 1.22762f
C456 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_10 VSS 1.22562f
C457 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_9 VSS 1.22562f
C458 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_8 VSS 1.22629f
C459 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_7 VSS 1.22696f
C460 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_6 VSS 1.22562f
C461 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_5 VSS 1.22562f
C462 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_4 VSS 1.22562f
C463 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_3 VSS 1.22629f
C464 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_2 VSS 1.22896f
C465 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_1 VSS 1.22562f
C466 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_0 VSS 1.22562f
C467 iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_2.di_tg_ctrl VSS 14.3155f
C468 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF6_0.vin VSS 4.48926f
C469 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inv_cross VSS 7.66312f
C470 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.buf_cross VSS 7.89561f
C471 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_1.inverter_NF2_1.vin VSS 2.82434f
C472 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS 3.36642f
C473 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS 3.36642f
C474 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VSS 2.49069f
C475 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS 3.36642f
C476 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS 3.36642f
C477 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS 3.36642f
C478 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS 3.36642f
C479 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS 3.36642f
C480 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0.S1 VSS 2.49069f
C481 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS 3.36642f
C482 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__nfet_01v8_lvt_WHJEU4_0.S1 VSS 3.36642f
C483 iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl_n VSS 11.5086f
C484 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_1.vin VSS 4.48926f
C485 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.transmission_gate_wo_dummy_0.v_b VSS 2.83622f
C486 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VSS 7.84314f
C487 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_7.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VSS 7.84314f
C488 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_1.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VSS 5.82216f
C489 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VSS 7.84314f
C490 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_8.vout VSS 51.5669f
C491 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_5.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VSS 7.84314f
C492 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_4.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VSS 7.84314f
C493 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutp VSS 74.2324f
C494 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_3.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VSS 7.84314f
C495 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_2.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VSS 7.84314f
C496 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF4_0.sky130_fd_pr__pfet_01v8_lvt_P4JB26_0.S1 VSS 5.82216f
C497 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_1.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VSS 7.84314f
C498 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_n_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_99 VSS 36.4777f
C499 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_6.vout VSS 75.0436f
C500 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.inverter_lv_en_NF6_0.sky130_fd_pr__pfet_01v8_lvt_P4QH36_0.S1 VSS 7.84314f
C501 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.ota_core_hybrid_bm_0.ota_core_en_n VSS 37.237f
C502 iq_modulator_half_0.passive_voltage_mode_mixer_0.transmission_gate_w_dummy_0.di_tg_ctrl VSS 14.3155f
C503 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF6_0.vin VSS 4.48926f
C504 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inv_cross VSS 7.66312f
C505 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.buf_cross VSS 7.89561f
C506 iq_modulator_half_0.passive_voltage_mode_mixer_0.lo_logic_0.inverter_NF2_1.vin VSS 2.82434f
C507 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.voutn VSS 74.9539f
C508 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_136 VSS 1.22562f
C509 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_135 VSS 1.22562f
C510 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_134 VSS 1.22562f
C511 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_133 VSS 1.22562f
C512 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_132 VSS 1.22696f
C513 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_131 VSS 1.22562f
C514 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_130 VSS 1.22562f
C515 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_129 VSS 1.22562f
C516 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_128 VSS 1.22629f
C517 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_127 VSS 1.22562f
C518 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_126 VSS 1.22562f
C519 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_125 VSS 1.22562f
C520 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_124 VSS 1.22562f
C521 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_123 VSS 1.22629f
C522 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_122 VSS 1.22696f
C523 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_121 VSS 1.22562f
C524 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_120 VSS 1.22562f
C525 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_119 VSS 1.22629f
C526 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_118 VSS 1.22629f
C527 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_117 VSS 1.22562f
C528 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_116 VSS 1.22562f
C529 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_115 VSS 1.22562f
C530 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_114 VSS 1.22562f
C531 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_113 VSS 1.22562f
C532 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_112 VSS 1.22696f
C533 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_111 VSS 1.22562f
C534 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_110 VSS 1.22562f
C535 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_109 VSS 1.22562f
C536 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_108 VSS 1.22629f
C537 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_107 VSS 1.22696f
C538 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_106 VSS 1.22562f
C539 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_105 VSS 1.22562f
C540 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_104 VSS 1.22562f
C541 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_103 VSS 1.22629f
C542 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_102 VSS 1.22696f
C543 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_101 VSS 1.22562f
C544 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_100 VSS 1.22562f
C545 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_99 VSS 36.1864f
C546 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_98 VSS 1.22629f
C547 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_97 VSS 1.22562f
C548 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_96 VSS 1.22562f
C549 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_95 VSS 1.22562f
C550 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_94 VSS 1.22562f
C551 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_93 VSS 1.22629f
C552 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_92 VSS 1.22696f
C553 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_91 VSS 1.22562f
C554 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_90 VSS 1.22562f
C555 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_89 VSS 1.22629f
C556 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_88 VSS 1.22629f
C557 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_87 VSS 1.22562f
C558 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_86 VSS 1.22562f
C559 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_85 VSS 1.22562f
C560 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_84 VSS 1.22562f
C561 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_83 VSS 1.22629f
C562 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_82 VSS 1.22696f
C563 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_81 VSS 1.22562f
C564 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_80 VSS 1.22562f
C565 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_79 VSS 1.22562f
C566 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_78 VSS 1.22629f
C567 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_77 VSS 1.22562f
C568 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_76 VSS 1.22562f
C569 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_75 VSS 1.22562f
C570 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_74 VSS 1.22562f
C571 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_73 VSS 1.22629f
C572 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_72 VSS 1.22562f
C573 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_71 VSS 1.22562f
C574 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_70 VSS 1.22562f
C575 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_69 VSS 1.22562f
C576 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_68 VSS 1.22629f
C577 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_67 VSS 1.22696f
C578 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_66 VSS 1.22562f
C579 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_65 VSS 1.22562f
C580 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_64 VSS 1.22562f
C581 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_63 VSS 1.22629f
C582 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_62 VSS 1.22696f
C583 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_61 VSS 1.22562f
C584 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_60 VSS 1.22562f
C585 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_59 VSS 1.22562f
C586 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_58 VSS 1.22562f
C587 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_57 VSS 1.22696f
C588 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_56 VSS 1.22562f
C589 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_55 VSS 1.22562f
C590 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_54 VSS 1.22562f
C591 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_53 VSS 1.22629f
C592 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_52 VSS 1.22696f
C593 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_51 VSS 1.22562f
C594 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_50 VSS 1.22562f
C595 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_49 VSS 1.22562f
C596 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_48 VSS 1.22629f
C597 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_47 VSS 1.22562f
C598 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_46 VSS 1.22562f
C599 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_45 VSS 1.22562f
C600 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_44 VSS 1.22562f
C601 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_43 VSS 1.22629f
C602 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_42 VSS 1.22696f
C603 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_41 VSS 1.22562f
C604 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_40 VSS 1.22562f
C605 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_39 VSS 1.22562f
C606 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_38 VSS 1.22629f
C607 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_37 VSS 1.22562f
C608 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC2p VSS 56.026f
C609 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_35 VSS 1.22562f
C610 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_34 VSS 1.22562f
C611 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_33 VSS 1.22629f
C612 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_32 VSS 1.22696f
C613 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_31 VSS 1.22562f
C614 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_30 VSS 1.22562f
C615 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_29 VSS 1.22562f
C616 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_28 VSS 1.22629f
C617 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_27 VSS 1.22562f
C618 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_26 VSS 1.22562f
C619 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_25 VSS 1.22562f
C620 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_24 VSS 1.22562f
C621 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_23 VSS 1.22629f
C622 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_22 VSS 1.22696f
C623 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_21 VSS 1.22562f
C624 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_20 VSS 1.22562f
C625 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_19 VSS 1.22562f
C626 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_18 VSS 1.22629f
C627 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.vC1p VSS 78.8372f
C628 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_16 VSS 1.22562f
C629 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_15 VSS 1.22562f
C630 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_14 VSS 1.22562f
C631 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_13 VSS 1.22562f
C632 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_12 VSS 1.22696f
C633 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_11 VSS 1.22562f
C634 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_10 VSS 1.22562f
C635 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_9 VSS 1.22562f
C636 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_8 VSS 1.22629f
C637 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_7 VSS 1.22562f
C638 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_6 VSS 1.22562f
C639 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_5 VSS 1.22562f
C640 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_4 VSS 1.22562f
C641 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_3 VSS 1.22896f
C642 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_2 VSS 1.22562f
C643 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R2_1 VSS 1.22562f
C644 iq_modulator_half_0.third_order_mfb_lp_filter_wo_C_0.resistors_0/resistors_p_0/sky130_fd_pr__res_xhigh_po_0p35_6YX8Z4_0.R1_0 VSS 1.22562f
.ends

