magic
tech sky130A
magscale 1 2
timestamp 1762641840
<< locali >>
rect -130 4680 1755 4695
rect -130 4550 -115 4680
rect 1740 4550 1755 4680
rect -130 4365 325 4550
rect 1295 4365 1755 4550
rect -130 4230 1755 4365
rect -130 4065 20 4230
rect -130 2290 -100 4065
rect -60 2290 20 4065
rect -130 2155 20 2290
rect 1600 4065 1755 4230
rect 1600 2290 1680 4065
rect 1720 2290 1755 4065
rect 1600 2155 1755 2290
rect -130 2130 1755 2155
rect -130 2095 20 2130
rect 1600 2095 1755 2130
rect -130 1925 1755 1985
rect -130 1800 20 1925
rect -130 1220 -100 1800
rect -60 1220 20 1800
rect -130 1070 20 1220
rect 1600 1800 1755 1925
rect 1600 1220 1680 1800
rect 1720 1220 1755 1800
rect 1600 1070 1755 1220
rect -130 925 1755 1070
rect -130 740 325 925
rect 1295 740 1755 925
rect -130 620 -115 740
rect 1740 620 1755 740
rect -130 605 1755 620
<< viali >>
rect -115 4550 1740 4680
rect 325 4365 1295 4550
rect -100 2290 -60 4065
rect 1680 2290 1720 4065
rect -100 1220 -60 1800
rect 1680 1220 1720 1800
rect 325 740 1295 925
rect -115 620 1740 740
<< metal1 >>
rect -130 4680 1755 4695
rect -130 4550 -115 4680
rect 1740 4550 1755 4680
rect -130 4535 325 4550
rect -130 4080 15 4535
rect 70 4435 240 4450
rect 70 4315 85 4435
rect 225 4315 240 4435
rect 310 4365 325 4535
rect 1295 4535 1755 4550
rect 1295 4365 1310 4535
rect 310 4350 1310 4365
rect 1370 4435 1540 4450
rect 70 4130 240 4315
rect 1370 4315 1385 4435
rect 1525 4315 1540 4435
rect 290 4135 1330 4295
rect 290 4080 375 4135
rect -130 4065 235 4080
rect -130 2290 -100 4065
rect -60 2290 85 4065
rect 225 2290 235 4065
rect -130 2275 235 2290
rect 270 2275 375 4080
rect 475 4070 635 4080
rect 475 2285 485 4070
rect 625 2285 635 4070
rect 475 2275 635 2285
rect 730 2275 890 4135
rect 1245 4080 1330 4135
rect 1370 4130 1540 4315
rect 1595 4080 1755 4535
rect 985 4070 1145 4080
rect 985 2285 995 4070
rect 1135 2285 1145 4070
rect 985 2275 1145 2285
rect 1245 2275 1405 4080
rect 1570 4065 1755 4080
rect 1570 2290 1680 4065
rect 1720 2290 1755 4065
rect 1570 2280 1755 2290
rect 1565 2275 1755 2280
rect 330 2195 1300 2230
rect -165 1885 1300 2195
rect 330 1850 1300 1885
rect -130 1800 55 1810
rect -130 1220 -100 1800
rect -60 1220 55 1800
rect -130 1215 55 1220
rect -130 1205 60 1215
rect 215 1210 375 1810
rect 475 1800 635 1810
rect 475 1220 485 1800
rect 625 1220 635 1800
rect 475 1210 635 1220
rect -130 755 15 1205
rect 70 985 240 1170
rect 290 1155 375 1210
rect 730 1155 890 1810
rect 985 1800 1145 1810
rect 985 1220 995 1800
rect 1135 1220 1145 1800
rect 985 1210 1145 1220
rect 1245 1210 1405 1810
rect 1570 1800 1755 1810
rect 1570 1220 1680 1800
rect 1720 1220 1755 1800
rect 1570 1215 1755 1220
rect 1245 1155 1330 1210
rect 1565 1205 1755 1215
rect 290 995 1330 1155
rect 70 865 85 985
rect 225 865 240 985
rect 1370 985 1540 1170
rect 70 850 240 865
rect 310 925 1310 940
rect 310 755 325 925
rect -130 740 325 755
rect 1295 755 1310 925
rect 1370 865 1385 985
rect 1525 865 1540 985
rect 1370 850 1540 865
rect 1595 755 1755 1205
rect 1295 740 1755 755
rect -130 620 -115 740
rect 1740 620 1755 740
rect -130 605 1755 620
<< via1 >>
rect 85 4315 225 4435
rect 1385 4315 1525 4435
rect 85 2290 225 4065
rect 485 2285 625 4070
rect 995 2285 1135 4070
rect 485 1220 625 1800
rect 995 1220 1135 1800
rect 85 865 225 985
rect 1385 865 1525 985
<< metal2 >>
rect -165 4435 1540 4450
rect -165 4315 85 4435
rect 225 4315 1385 4435
rect 1525 4315 1540 4435
rect -165 4300 1540 4315
rect 70 4065 240 4080
rect 70 2290 85 4065
rect 225 2290 240 4065
rect 70 1000 240 2290
rect 475 4070 635 4080
rect 475 2285 485 4070
rect 625 2285 635 4070
rect 475 2240 635 2285
rect 985 4070 1145 4080
rect 985 2285 995 4070
rect 1135 2285 1145 4070
rect 985 2240 1145 2285
rect 475 1840 1770 2240
rect 475 1800 635 1840
rect 475 1220 485 1800
rect 625 1220 635 1800
rect 475 1210 635 1220
rect 985 1800 1145 1840
rect 985 1220 995 1800
rect 1135 1220 1145 1800
rect 985 1210 1145 1220
rect 70 985 1540 1000
rect 70 865 85 985
rect 225 865 1385 985
rect 1525 865 1540 985
rect 70 850 1540 865
use sky130_fd_pr__nfet_01v8_lvt_XCBGUP  sky130_fd_pr__nfet_01v8_lvt_XCBGUP_0
timestamp 1762641840
transform 1 0 811 0 1 1510
box -941 -510 941 510
use sky130_fd_pr__pfet_01v8_lvt_P4JB26  sky130_fd_pr__pfet_01v8_lvt_P4JB26_0
timestamp 1762641840
transform 1 0 811 0 1 3179
box -941 -1119 941 1119
<< labels >>
flabel metal2 -155 4370 -155 4370 0 FreeSans 320 0 0 0 di_en
port 8 nsew
flabel viali 965 4610 965 4610 0 FreeSans 400 0 0 0 VDD
port 11 nsew
flabel metal1 -155 2040 -155 2040 0 FreeSans 320 0 0 0 vin
port 12 nsew
flabel metal2 1760 2040 1760 2040 0 FreeSans 320 0 0 0 vout
port 14 nsew
flabel viali 1040 670 1040 670 0 FreeSans 400 0 0 0 VSS
port 10 nsew
<< end >>
